RC Circuit Transient Response
****** Discrete Bipolar Electrical Parameters ******
** NPN Epitaxial Silicon Transistor
** Package: D-PAK / TO-220
** High Voltage Power Switching Application
**---------------------------------------------------------------------------
.SUBCKT KSC5502D C B E
q1 C B E VNPN
d1 E C   DFW

.MODEL VNPN npn (                               
+ IS = 1.4547E-12      BF = 58.7             NF = 1               
+ BR = 20.4            NR = 1                ISE = 2.8201E-10     
+ NE = 2.0             ISC = 2.2481E-7       NC = 1.5              
+ VAF = 18             VAR = 100             IKF = 0.1246           
+ IKR = 0.06           RB = 2.83             RBM = 0.0631          
+ IRB = 0.000210       RE = 0.02             RC = 0.04             
+ CJE = 8.2308E-10     VJE = 0.6678          MJE = 0.3289          
+ FC = 0.5             CJC = 1.9684E-10      VJC = 0.4527
+ MJC = 0.6368         XTB = 1.1034          EG = 0.95
+ XTI = 3              TF = 1.4076E-8  )

.MODEL DFW d (
+ IS = 2.4E-13         N = 1                 RS = 0.052   
+ EG = 1.158           CJO = 1E-10 )
.ENDS
**---------------------------------------------------------------------------
** Creation: Sep.-26-2007
** Fairchild Semiconductor




*****************************************************************
* INFINEON Power Transistors                                    *
* Level-1 / 3 PSPICE Library for small signal transistors       *
* Version 270715                                                *
*                                                               *
*                                                               *
* Models provided by Infineon are not warranted by Infineon as  *
* fully representing all the specifications and operating       *
* characteristics of the semiconductor product to which the     *
* model relates. The models describe the characteristics of     *
* typical devices.                                              *
* In all cases, the current data sheet information for a given  *
* device is the final design guideline and the only actual      *
* performance specification.                                    *
* Although models can be a useful tool in evaluating device     *
* performance, they cannot model exact device performance under *
* all conditions, nor are they intended to replace bread-       *
* boarding for final verification. INFINEON therefore does not  *
* assume any liability arising from their use.                  *
* INFINEON reserves the right to change models without prior    *
* notice.                                                       *
*                                                               *
*****************************************************************
*                                                               *
*   BSS131         (n-channel, 240 V enhancement)               *
*   BSS87          (n-channel, 240 V enhancement)               *
*   BSP89          (n-channel, 240 V enhancement)               *
*   BSP88          (n-channel, 240 V enhancement)               *
*   BSP129         (n-channel, 240 V depletion)                 *
*   SISC0_97N24D   (n-channel, 240 V depletion)                 *
*   BSS139         (n-channel, 250 V depletion)                 *
*   BSP324         (n-channel, 400 V enhancement)               *
*   SISC1_4N40E    (n-channel, 400 V enhancement                *   
*   BSP125         (n-channel, 600 V enhancement)               *
*   BSS225         (n-channel, 600 V enhancement)               *
*   BSS127         (n-channel, 600 V enhancement)               *
*   BSP135         (n-channel, 600 V depletion)                 *
*   SISC1_4N60D    (n-channel, 600 V depletion)                 *
*   BSS126         (n-channel, 600 V depletion)                 *
*   BSP300         (n-channel, 800 V enhancement, Level 0 only) *
*                                                               *
*****************************************************************
* thermal nodes of level 3 models:                              *
*                                                               *
*  .SUBCKT BSP135 drain gate source Tj Tcase                    *
*  Tj :    potential=temperature (in °C) at junction (typically *
*          not connected)                                       *
*  Tcase/Tsolder_joint :                                        *
*          node where the boundary contition - external heat    *
*          sinks etc - have to be connected (ideal heat sink    *
*          can be modeled by using a voltage source stating the *
*          ambient temperature in °C between Tcase and ground.  *
*                                                               *  
*****************************************************************
   
 

.SUBCKT K_240_a_var dd g s Tj PARAMS: a=1 dVth=0 dR=0 dgfs=0 Inn=1 Unn=1 Rmax=1
+gmin=1 Rs=1 Rp=1 dC=0 heat=1

.PARAM  Vth0=1.45      beta4c=0.217   ph0=25.7       ph1=0.038      Ubr=290
.PARAM  Rd=1.95        nmu=2.6        Rf=0.2         rpa=0.06877    lnIsj=-24.7
.PARAM  Rdi=0.2

.PARAM  Tref=298     T0=273      auth=3m      c=0.82       mu_bet=0.4
.PARAM  f_bet=-2     ndi=1.2     UTnbr=207m   lnBr=-23     kbq=85.8u
.PARAM  Wcml={beta4c*4*c}        
.PARAM  aubr={0.93m*UBr}
.PARAM  dvgs={0.1-0.06*Vth0}

.PARAM  f1=65p         f2=92p         f3=198p        f4=265p        f5=290p
.PARAM  U0=0.5         nd=0.44        nc=0.5         g1=1.9         bb=-3
.PARAM  sl=65p         remp=0p        ta=60n         td=20n

.PARAM  Vmin=0.8       Vmax=1.8       dCmax=0.35
.PARAM  Vth={Vth0+(Vmax-Vth0)*limit(dVth,0,1)-(Vmin-Vth0)*limit(dVth,-1,0)}
.PARAM  p0={Wcml*a*((1-f_bet)*(T0/Tref)**mu_bet+f_bet)    }
.PARAM  Rlim={(Rmax-Rs-(Unn-Vth0-Inn*Rs-SQRT((Unn-Vth0-Inn*Rs)**2-4*c*Inn/p0))/(2*c*Inn))/(1+rpa*(Inn/a)**2)} 
.PARAM  dRd={Rd/a+if(dVth==0,limit(dR,0,1)*max(Rlim-Rd/a,0),0)} 
.PARAM  bet={Wcml}

.PARAM  dC1={1+dCmax*limit(dC,0,1)} 
.PARAM  Cox={f1*a*dC1}
.PARAM  Cds0={f2*a*dC1}
.PARAM  Cgs0={f3*a*dC1}
.PARAM  Cox1={f5*a*dC1}
.PARAM  Crand={remp*SQRT(a)}
.PARAM  dRdi={Rdi/a}

.FUNC U1(Uds,T)       {(SQRT(1+4*(0.4+(T-T0-25)*2m)*abs(Uds))-1)/2/(0.4+(T-T0-25)*2m)}
.FUNC I2(p,Uee,z1,pp) {if(Uee>pp,(Uee-c*z1)*z1,p*(pp-p)/c*exp((Uee-pp-(min(0,Uee))**2)/p))}
.FUNC Ig(Uds,T,p,Uee) {bet*((1-f_bet)*(T0/T)**mu_bet+f_bet)*I2(p,Uee,min(Uds,Uee/(2*c)),min(2*p,p+c*Uds))}
.FUNC Iges(Uds,Ugs,T) 
 +{a*(sgn(Uds)*Ig(U1(Uds,T),T,1/(ph0-ph1*T),Ugs-Vth+auth*(T-Tref))+exp(min(lnBr+(abs(Uds)-UBr-aubr*(T-Tref))/UTnbr,25)))}

.FUNC Isjt(Tj)           {exp(min(lnIsj+(Tj/Tref-1)*1.12/(ndi*kbq*Tj),9))*(Tj/Tref)**1.5}
.FUNC Idiode(Usd,Tj,Iss) {exp(min(log(Iss)+Usd/(ndi*kbq*Tj),9))-Iss}
.FUNC Idiod(Usd,Tj)      {a*Idiode(Usd,Tj,Isjt(Tj))}

.FUNC QCdg(x,z)  {if(f4>f5,(f5**2-(f4-z*sl)**2)/(2*sl)+f5*min(x,(f4-f5)/sl),f4*z-sl*z**2/2-f5*max((f4-f5)/sl-x,0))}

E_Edg     d   ox  VALUE {V(d,g)-(min(V(d,g),-bb)+1/(g1*(1-nc))*((1/(1+g1*max(V(d,g)+bb,0)))**(nc-1)-1))}
C_Cdg     ox  g   {Cox}
E_Edg1    d   ox1 VALUE {V(d,g)-QCdg(V(d,g),limit(V(d,g),(f4-f5)/sl,f4/sl))/f5}
C_Cdg1    ox1 g   {Cox1}
C_Cdg2    d   g   {Crand}

E_Eds     d edep  VALUE {(V(d2,s)-I(V_sense3)/Cds0)}
C_Cds  edep    s  {Cds0}
C_Cds2   d2    s  {Cds0/500}

C_Cgs     g    s  {Cgs0}

G_chan    d    s  VALUE={Iges(V(d,s),V(g,s),T0+limit(V(Tj),-200,350))}
E_RMos   d1    d  VALUE={I(V_sense)*(Rf*dRd+(1-Rf)*dRd*((limit(V(Tj),-200,999)+T0)/Tref)**nmu)*(1+rpa*(I(V_sense)/a)**2)}
V_sense  dd   d1  0
G_diode   s   d2  VALUE={Idiod(V(s,d2),T0+limit(V(Tj),-200,499))}
R_Rdio   d2   d3  {dRdi}
V_sense2 d1   d3  0

L_L001    a    c  {td/(ta+td)}
R_R001    a    b  {1/ta}
V_sense3  c    f  0
R_sense3  f    0  1
E_E001    b    0  VALUE {I(V_sense2)}
E_E002    e    0  VALUE {1Meg*Cds0*(1/(1-nd)*U0**nd*(limit(U0+V(d2,s),U0/2,2*UBr))**(1-nd)+2**nd*min(V(d2,s)+U0/2,0))}
R_R002    e    c  1Meg

R1        g    s  1G
Rd01      d    s  500Meg
Rd02     d2    s  500Meg
Rd03     d1    d  10k

G_TH      0    Tj  VALUE = {heat*LIMIT(I(V_sense)*V(dd,s),0,100k)}

.ENDS
*$

**************************************************************************************


.SUBCKT K_240_b_var dd g s Tj PARAMS: a=1 dVth=0 dR=0 dgfs=0 Inn=1 Unn=1 Rmax=1
+gmin=1 Rs=1 Rp=1 dC=0 heat=1

.PARAM  Vth0=1.5       beta4c=0.243   ph0=25.7       ph1=0.038      Ubr=290
.PARAM  Rd=1.95        nmu=2.6        Rf=0.2         rpa=0.06877    lnIsj=-24.7
.PARAM  Rdi=0.2

.PARAM  Tref=298     T0=273      auth=3m      c=0.82       mu_bet=0.4
.PARAM  f_bet=-2     ndi=1.2     UTnbr=207m   lnBr=-23     kbq=85.8u
.PARAM  Wcml={beta4c*4*c}        
.PARAM  aubr={0.93m*UBr}
.PARAM  dvgs={0.1-0.06*Vth0}

.PARAM  f1=65p         f2=69p         f3=139p        f4=310p        f5=270p
.PARAM  U0=0.5         nd=0.47        nc=0.5         g1=1.9         bb=-3.3
.PARAM  sl=65p         remp=0p        ta=60n         td=20n

.PARAM  Vmin=0.8       Vmax=1.8       dCmax=0.35
.PARAM  Vth={Vth0+(Vmax-Vth0)*limit(dVth,0,1)-(Vmin-Vth0)*limit(dVth,-1,0)}
.PARAM  p0={Wcml*a*((1-f_bet)*(T0/Tref)**mu_bet+f_bet)    }
.PARAM  Rlim={(Rmax-Rs-(Unn-Vth0-Inn*Rs-SQRT((Unn-Vth0-Inn*Rs)**2-4*c*Inn/p0))/(2*c*Inn))/(1+rpa*(Inn/a)**2)} 
.PARAM  dRd={Rd/a+if(dVth==0,limit(dR,0,1)*max(Rlim-Rd/a,0),0)} 
.PARAM  bet={Wcml}

.PARAM  dC1={1+dCmax*limit(dC,0,1)} 
.PARAM  Cox={f1*a*dC1}
.PARAM  Cds0={f2*a*dC1}
.PARAM  Cgs0={f3*a*dC1}
.PARAM  Cox1={f5*a*dC1}
.PARAM  Crand={remp*SQRT(a)}
.PARAM  dRdi={Rdi/a}

.FUNC U1(Uds,T)       {(SQRT(1+4*(0.4+(T-T0-25)*2m)*abs(Uds))-1)/2/(0.4+(T-T0-25)*2m)}
.FUNC I2(p,Uee,z1,pp) {if(Uee>pp,(Uee-c*z1)*z1,p*(pp-p)/c*exp((Uee-pp-(min(0,Uee))**2)/p))}
.FUNC Ig(Uds,T,p,Uee) {bet*((1-f_bet)*(T0/T)**mu_bet+f_bet)*I2(p,Uee,min(Uds,Uee/(2*c)),min(2*p,p+c*Uds))}
.FUNC Iges(Uds,Ugs,T) 
 +{a*(sgn(Uds)*Ig(U1(Uds,T),T,1/(ph0-ph1*T),Ugs-Vth+auth*(T-Tref))+exp(min(lnBr+(abs(Uds)-UBr-aubr*(T-Tref))/UTnbr,25)))}

.FUNC Isjt(Tj)           {exp(min(lnIsj+(Tj/Tref-1)*1.12/(ndi*kbq*Tj),9))*(Tj/Tref)**1.5}
.FUNC Idiode(Usd,Tj,Iss) {exp(min(log(Iss)+Usd/(ndi*kbq*Tj),9))-Iss}
.FUNC Idiod(Usd,Tj)      {a*Idiode(Usd,Tj,Isjt(Tj))}

.FUNC QCdg(x,z)  {if(f4>f5,(f5**2-(f4-z*sl)**2)/(2*sl)+f5*min(x,(f4-f5)/sl),f4*z-sl*z**2/2-f5*max((f4-f5)/sl-x,0))}

E_Edg     d   ox  VALUE {V(d,g)-(min(V(d,g),-bb)+1/(g1*(1-nc))*((1/(1+g1*max(V(d,g)+bb,0)))**(nc-1)-1))}
C_Cdg     ox  g   {Cox}
E_Edg1    d   ox1 VALUE {V(d,g)-QCdg(V(d,g),limit(V(d,g),(f4-f5)/sl,f4/sl))/f5}
C_Cdg1    ox1 g   {Cox1}
C_Cdg2    d   g   {Crand}

E_Eds     d edep  VALUE {(V(d2,s)-I(V_sense3)/Cds0)}
C_Cds  edep    s  {Cds0}
C_Cds2   d2    s  {Cds0/500}

C_Cgs     g    s  {Cgs0}

G_chan    d    s  VALUE={Iges(V(d,s),V(g,s),T0+limit(V(Tj),-200,350))}
E_RMos   d1    d  VALUE={I(V_sense)*(Rf*dRd+(1-Rf)*dRd*((limit(V(Tj),-200,999)+T0)/Tref)**nmu)*(1+rpa*(I(V_sense)/a)**2)}
V_sense  dd   d1  0
G_diode   s   d2  VALUE={Idiod(V(s,d2),T0+limit(V(Tj),-200,499))}
R_Rdio   d2   d3  {dRdi}
V_sense2 d1   d3  0

L_L001    a    c  {td/(ta+td)}
R_R001    a    b  {1/ta}
V_sense3  c    f  0
R_sense3  f    0  1
E_E001    b    0  VALUE {I(V_sense2)}
E_E002    e    0  VALUE {1Meg*Cds0*(1/(1-nd)*U0**nd*(limit(U0+V(d2,s),U0/2,2*UBr))**(1-nd)+2**nd*min(V(d2,s)+U0/2,0))}
R_R002    e    c  1Meg

R1        g    s  1G
Rd01      d    s  500Meg
Rd02     d2    s  500Meg
Rd03     d1    d  10k

G_TH      0    Tj  VALUE = {heat*LIMIT(I(V_sense)*V(dd,s),0,100k)}

.ENDS
*$

**************************************************************************************


.SUBCKT K_240_c_var dd g s Tj PARAMS: a=1 dVth=0 dR=0 dgfs=0 Inn=1 Unn=1 Rmax=1
+gmin=1 Rs=1 Rp=1 dC=0 heat=1

.PARAM  Vth0=1.1       beta4c=0.243   ph0=25.7       ph1=0.038      Ubr=290
.PARAM  Rd=1.95        nmu=2.6        Rf=0.2         rpa=0.06877    lnIsj=-24.7
.PARAM  Rdi=0.2

.PARAM  Tref=298     T0=273      auth=3m      c=0.82       mu_bet=0.4
.PARAM  f_bet=-2     ndi=1.2     UTnbr=207m   lnBr=-23     kbq=85.8u
.PARAM  Wcml={beta4c*4*c}        
.PARAM  aubr={0.93m*UBr}
.PARAM  dvgs={0.1-0.06*Vth0}

.PARAM  f1=65p         f2=69p         f3=139p        f4=310p        f5=270p
.PARAM  U0=0.5         nd=0.47        nc=0.5         g1=1.9         bb=-3.3
.PARAM  sl=65p         remp=0p        ta=60n         td=20n

.PARAM  Vmin=0.6       Vmax=1.4       dCmax=0.35
.PARAM  Vth={Vth0+(Vmax-Vth0)*limit(dVth,0,1)-(Vmin-Vth0)*limit(dVth,-1,0)}
.PARAM  p0={Wcml*a*((1-f_bet)*(T0/Tref)**mu_bet+f_bet)    }
.PARAM  Rlim={(Rmax-Rs-(Unn-Vth0-Inn*Rs-SQRT((Unn-Vth0-Inn*Rs)**2-4*c*Inn/p0))/(2*c*Inn))/(1+rpa*(Inn/a)**2)} 
.PARAM  dRd={Rd/a+if(dVth==0,limit(dR,0,1)*max(Rlim-Rd/a,0),0)} 
.PARAM  bet={Wcml}

.PARAM  dC1={1+dCmax*limit(dC,0,1)} 
.PARAM  Cox={f1*a*dC1}
.PARAM  Cds0={f2*a*dC1}
.PARAM  Cgs0={f3*a*dC1}
.PARAM  Cox1={f5*a*dC1}
.PARAM  Crand={remp*SQRT(a)}
.PARAM  dRdi={Rdi/a}

.FUNC U1(Uds,T)       {(SQRT(1+4*(0.4+(T-T0-25)*2m)*abs(Uds))-1)/2/(0.4+(T-T0-25)*2m)}
.FUNC I2(p,Uee,z1,pp) {if(Uee>pp,(Uee-c*z1)*z1,p*(pp-p)/c*exp((Uee-pp-(min(0,Uee))**2)/p))}
.FUNC Ig(Uds,T,p,Uee) {bet*((1-f_bet)*(T0/T)**mu_bet+f_bet)*I2(p,Uee,min(Uds,Uee/(2*c)),min(2*p,p+c*Uds))}
.FUNC Iges(Uds,Ugs,T) 
 +{a*(sgn(Uds)*Ig(U1(Uds,T),T,1/(ph0-ph1*T),Ugs-Vth+auth*(T-Tref))+exp(min(lnBr+(abs(Uds)-UBr-aubr*(T-Tref))/UTnbr,25)))}

.FUNC Isjt(Tj)           {exp(min(lnIsj+(Tj/Tref-1)*1.12/(ndi*kbq*Tj),9))*(Tj/Tref)**1.5}
.FUNC Idiode(Usd,Tj,Iss) {exp(min(log(Iss)+Usd/(ndi*kbq*Tj),9))-Iss}
.FUNC Idiod(Usd,Tj)      {a*Idiode(Usd,Tj,Isjt(Tj))}

.FUNC QCdg(x,z)  {if(f4>f5,(f5**2-(f4-z*sl)**2)/(2*sl)+f5*min(x,(f4-f5)/sl),f4*z-sl*z**2/2-f5*max((f4-f5)/sl-x,0))}

E_Edg     d   ox  VALUE {V(d,g)-(min(V(d,g),-bb)+1/(g1*(1-nc))*((1/(1+g1*max(V(d,g)+bb,0)))**(nc-1)-1))}
C_Cdg     ox  g   {Cox}
E_Edg1    d   ox1 VALUE {V(d,g)-QCdg(V(d,g),limit(V(d,g),(f4-f5)/sl,f4/sl))/f5}
C_Cdg1    ox1 g   {Cox1}
C_Cdg2    d   g   {Crand}

E_Eds     d edep  VALUE {(V(d2,s)-I(V_sense3)/Cds0)}
C_Cds  edep    s  {Cds0}
C_Cds2   d2    s  {Cds0/500}

C_Cgs     g    s  {Cgs0}

G_chan    d    s  VALUE={Iges(V(d,s),V(g,s),T0+limit(V(Tj),-200,350))}
E_RMos   d1    d  VALUE={I(V_sense)*(Rf*dRd+(1-Rf)*dRd*((limit(V(Tj),-200,999)+T0)/Tref)**nmu)*(1+rpa*(I(V_sense)/a)**2)}
V_sense  dd   d1  0
G_diode   s   d2  VALUE={Idiod(V(s,d2),T0+limit(V(Tj),-200,499))}
R_Rdio   d2   d3  {dRdi}
V_sense2 d1   d3  0

L_L001    a    c  {td/(ta+td)}
R_R001    a    b  {1/ta}
V_sense3  c    f  0
R_sense3  f    0  1
E_E001    b    0  VALUE {I(V_sense2)}
E_E002    e    0  VALUE {1Meg*Cds0*(1/(1-nd)*U0**nd*(limit(U0+V(d2,s),U0/2,2*UBr))**(1-nd)+2**nd*min(V(d2,s)+U0/2,0))}
R_R002    e    c  1Meg

R1        g    s  1G
Rd01      d    s  500Meg
Rd02     d2    s  500Meg
Rd03     d1    d  10k

G_TH      0    Tj  VALUE = {heat*LIMIT(I(V_sense)*V(dd,s),0,100k)}

.ENDS
*$

**************************************************************************************


.SUBCKT K_240_d_var dd g s Tj PARAMS: a=1 dVth=0 dR=0 dgfs=0 Inn=1 Unn=1 Rmax=1
+gmin=1 Rs=1 Rp=1 dC=0 heat=1

.PARAM  Vth0=-1.05     beta4c=0.243   ph0=20         ph1=0.026      Ubr=290
.PARAM  Rd=1.95        nmu=2.6        Rf=0.2         rpa=0.06877    lnIsj=-24.7
.PARAM  Rdi=0.2

.PARAM  Tref=298     T0=273      auth=3m      c=0.82       mu_bet=0.4
.PARAM  f_bet=-2     ndi=1.2     UTnbr=207m   lnBr=-23     kbq=85.8u
.PARAM  Wcml={beta4c*4*c}        
.PARAM  aubr={0.93m*UBr}
.PARAM  dvgs={0.1-0.06*Vth0}

.PARAM  f1=65p         f2=69p         f3=139p        f4=360p        f5=270p
.PARAM  U0=0.5         nd=0.47        nc=0.5         g1=1.9         bb=-7
.PARAM  sl=45p         remp=0p        ta=60n         td=20n

.PARAM  Vmin=-1.75      Vmax=-0.65        dCmax=0.35
.PARAM  Vth={Vth0+(Vmax-Vth0)*limit(dVth,0,1)-(Vmin-Vth0)*limit(dVth,-1,0)}
.PARAM  p0={Wcml*a*((1-f_bet)*(T0/Tref)**mu_bet+f_bet)    }
.PARAM  Rlim={(Rmax-Rs-(Unn-Vth0-Inn*Rs-SQRT((Unn-Vth0-Inn*Rs)**2-4*c*Inn/p0))/(2*c*Inn))/(1+rpa*(Inn/a)**2)} 
.PARAM  dRd={Rd/a+if(dVth==0,limit(dR,0,1)*max(Rlim-Rd/a,0),0)} 
.PARAM  bet={Wcml}

.PARAM  dC1={1+dCmax*limit(dC,0,1)} 
.PARAM  Cox={f1*a*dC1}
.PARAM  Cds0={f2*a*dC1}
.PARAM  Cgs0={f3*a*dC1}
.PARAM  Cox1={f5*a*dC1}
.PARAM  Crand={remp*SQRT(a)}
.PARAM  dRdi={Rdi/a}

.FUNC U1(Uds,T)       {(SQRT(1+4*(0.4+(T-T0-25)*2m)*abs(Uds))-1)/2/(0.4+(T-T0-25)*2m)}
.FUNC I2(p,Uee,z1,pp) {if(Uee>pp,(Uee-c*z1)*z1,p*(pp-p)/c*exp((Uee-pp-(min(0,Uee))**2)/p))}
.FUNC Ig(Uds,T,p,Uee) {bet*((1-f_bet)*(T0/T)**mu_bet+f_bet)*I2(p,Uee,min(Uds,Uee/(2*c)),min(2*p,p+c*Uds))}
.FUNC Iges(Uds,Ugs,T) 
 +{a*(sgn(Uds)*Ig(U1(Uds,T),T,1/(ph0-ph1*T),Ugs-Vth+auth*(T-Tref))+exp(min(lnBr+(abs(Uds)-UBr-aubr*(T-Tref))/UTnbr,25)))}

.FUNC Isjt(Tj)           {exp(min(lnIsj+(Tj/Tref-1)*1.12/(ndi*kbq*Tj),9))*(Tj/Tref)**1.5}
.FUNC Idiode(Usd,Tj,Iss) {exp(min(log(Iss)+Usd/(ndi*kbq*Tj),9))-Iss}
.FUNC Idiod(Usd,Tj)      {a*Idiode(Usd,Tj,Isjt(Tj))}

.FUNC QCdg(x,z)  {if(f4>f5,(f5**2-(f4-z*sl)**2)/(2*sl)+f5*min(x,(f4-f5)/sl),f4*z-sl*z**2/2-f5*max((f4-f5)/sl-x,0))}

E_Edg     d   ox  VALUE {V(d,g)-(min(V(d,g),-bb)+1/(g1*(1-nc))*((1/(1+g1*max(V(d,g)+bb,0)))**(nc-1)-1))}
C_Cdg     ox  g   {Cox}
E_Edg1    d   ox1 VALUE {V(d,g)-QCdg(V(d,g),limit(V(d,g),(f4-f5)/sl,f4/sl))/f5}
C_Cdg1    ox1 g   {Cox1}
C_Cdg2    d   g   {Crand}

E_Eds     d edep  VALUE {(V(d2,s)-I(V_sense3)/Cds0)}
C_Cds  edep    s  {Cds0}
C_Cds2   d2    s  {Cds0/500}

C_Cgs     g    s  {Cgs0}

G_chan    d    s  VALUE={Iges(V(d,s),V(g,s),T0+limit(V(Tj),-200,350))}
E_RMos   d1    d  VALUE={I(V_sense)*(Rf*dRd+(1-Rf)*dRd*((limit(V(Tj),-200,999)+T0)/Tref)**nmu)*(1+rpa*(I(V_sense)/a)**2)}
V_sense  dd   d1  0
G_diode   s   d2  VALUE={Idiod(V(s,d2),T0+limit(V(Tj),-200,499))}
R_Rdio   d2   d3  {dRdi}
V_sense2 d1   d3  0

L_L001    a    c  {td/(ta+td)}
R_R001    a    b  {1/ta}
V_sense3  c    f  0
R_sense3  f    0  1
E_E001    b    0  VALUE {I(V_sense2)}
E_E002    e    0  VALUE {1Meg*Cds0*(1/(1-nd)*U0**nd*(limit(U0+V(d2,s),U0/2,2*UBr))**(1-nd)+2**nd*min(V(d2,s)+U0/2,0))}
R_R002    e    c  1Meg

R1        g    s  1G
Rd01      d    s  500Meg
Rd02     d2    s  500Meg
Rd03     d1    d  10k

G_TH      0    Tj  VALUE = {heat*LIMIT(I(V_sense)*V(dd,s),0,100k)}

.ENDS
*$

**************************************************************************************


.SUBCKT K_250_d_var dd g s Tj PARAMS: a=1 dVth=0 dR=0 dgfs=0 Inn=1 Unn=1 Rmax=1
+gmin=1 Rs=1 Rp=1 dC=0 heat=1

.PARAM  Vth0=-1.1      beta4c=0.217   ph0=20         ph1=0.026      Ubr=295
.PARAM  Rd=2           nmu=2.6        Rf=0.15        rpa=0.10933    lnIsj=-24.7
.PARAM  Rdi=0.2

.PARAM  Tref=298     T0=273      auth=3m      c=0.82       mu_bet=0.4
.PARAM  f_bet=-2     ndi=1.2     UTnbr=207m   lnBr=-23     kbq=85.8u
.PARAM  Wcml={beta4c*4*c}        
.PARAM  aubr={0.93m*UBr}
.PARAM  dvgs={0.1-0.06*Vth0}

.PARAM  f1=65p         f2=85p         f3=198p        f4=305p        f5=314p
.PARAM  U0=0.5         nd=0.45        nc=0.5         g1=2.2         bb=-7.5
.PARAM  sl=31p         remp=0p        ta=60n         td=20n

.PARAM  Vmin=-2.1      Vmax=-1        dCmax=0.35
.PARAM  Vth={Vth0+(Vmax-Vth0)*limit(dVth,0,1)-(Vmin-Vth0)*limit(dVth,-1,0)}
.PARAM  p0={Wcml*a*((1-f_bet)*(T0/Tref)**mu_bet+f_bet)    }
.PARAM  Rlim={(Rmax-Rs-(Unn-Vth0-Inn*Rs-SQRT((Unn-Vth0-Inn*Rs)**2-4*c*Inn/p0))/(2*c*Inn))/(1+rpa*(Inn/a)**2)} 
.PARAM  dRd={Rd/a+if(dVth==0,limit(dR,0,1)*max(Rlim-Rd/a,0),0)} 
.PARAM  bet={Wcml}

.PARAM  dC1={1+dCmax*limit(dC,0,1)} 
.PARAM  Cox={f1*a*dC1}
.PARAM  Cds0={f2*a*dC1}
.PARAM  Cgs0={f3*a*dC1}
.PARAM  Cox1={f5*a*dC1}
.PARAM  Crand={remp*SQRT(a)}
.PARAM  dRdi={Rdi/a}

.FUNC U1(Uds,T)       {(SQRT(1+4*(0.4+(T-T0-25)*2m)*abs(Uds))-1)/2/(0.4+(T-T0-25)*2m)}
.FUNC I2(p,Uee,z1,pp) {if(Uee>pp,(Uee-c*z1)*z1,p*(pp-p)/c*exp((Uee-pp-(min(0,Uee))**2)/p))}
.FUNC Ig(Uds,T,p,Uee) {bet*((1-f_bet)*(T0/T)**mu_bet+f_bet)*I2(p,Uee,min(Uds,Uee/(2*c)),min(2*p,p+c*Uds))}
.FUNC Iges(Uds,Ugs,T) 
 +{a*(sgn(Uds)*Ig(U1(Uds,T),T,1/(ph0-ph1*T),Ugs-Vth+auth*(T-Tref))+exp(min(lnBr+(abs(Uds)-UBr-aubr*(T-Tref))/UTnbr,25)))}

.FUNC Isjt(Tj)           {exp(min(lnIsj+(Tj/Tref-1)*1.12/(ndi*kbq*Tj),9))*(Tj/Tref)**1.5}
.FUNC Idiode(Usd,Tj,Iss) {exp(min(log(Iss)+Usd/(ndi*kbq*Tj),9))-Iss}
.FUNC Idiod(Usd,Tj)      {a*Idiode(Usd,Tj,Isjt(Tj))}

.FUNC QCdg(x,z)  {if(f4>f5,(f5**2-(f4-z*sl)**2)/(2*sl)+f5*min(x,(f4-f5)/sl),f4*z-sl*z**2/2-f5*max((f4-f5)/sl-x,0))}

E_Edg     d   ox  VALUE {V(d,g)-(min(V(d,g),-bb)+1/(g1*(1-nc))*((1/(1+g1*max(V(d,g)+bb,0)))**(nc-1)-1))}
C_Cdg     ox  g   {Cox}
E_Edg1    d   ox1 VALUE {V(d,g)-QCdg(V(d,g),limit(V(d,g),(f4-f5)/sl,f4/sl))/f5}
C_Cdg1    ox1 g   {Cox1}
C_Cdg2    d   g   {Crand}

E_Eds     d edep  VALUE {(V(d2,s)-I(V_sense3)/Cds0)}
C_Cds  edep    s  {Cds0}
C_Cds2   d2    s  {Cds0/500}

C_Cgs     g    s  {Cgs0}

G_chan    d    s  VALUE={Iges(V(d,s),V(g,s),T0+limit(V(Tj),-200,350))}
E_RMos   d1    d  VALUE={I(V_sense)*(Rf*dRd+(1-Rf)*dRd*((limit(V(Tj),-200,999)+T0)/Tref)**nmu)*(1+rpa*(I(V_sense)/a)**2)}
V_sense  dd   d1  0
G_diode   s   d2  VALUE={Idiod(V(s,d2),T0+limit(V(Tj),-200,499))}
R_Rdio   d2   d3  {dRdi}
V_sense2 d1   d3  0

L_L001    a    c  {td/(ta+td)}
R_R001    a    b  {1/ta}
V_sense3  c    f  0
R_sense3  f    0  1
E_E001    b    0  VALUE {I(V_sense2)}
E_E002    e    0  VALUE {1Meg*Cds0*(1/(1-nd)*U0**nd*(limit(U0+V(d2,s),U0/2,2*UBr))**(1-nd)+2**nd*min(V(d2,s)+U0/2,0))}
R_R002    e    c  1Meg

R1        g    s  1G
Rd01      d    s  500Meg
Rd02     d2    s  500Meg
Rd03     d1    d  10k

G_TH      0    Tj  VALUE = {heat*LIMIT(I(V_sense)*V(dd,s),0,100k)}

.ENDS
*$

**************************************************************************************


.SUBCKT K_400_a_var dd g s Tj PARAMS: a=1 dVth=0 dR=0 dgfs=0 Inn=1 Unn=1 Rmax=1
+gmin=1 Rs=1 Rp=1 dC=0 heat=1

.PARAM  Vth0=2.07      beta4c=0.157   ph0=25.7       ph1=0.038      Ubr=495
.PARAM  Rd=5.75        nmu=2.65       Rf=0.12        rpa=0.28717    lnIsj=-24.7
.PARAM  Rdi=0.2

.PARAM  Tref=298     T0=273      auth=3m      c=0.82       mu_bet=0.4
.PARAM  f_bet=-2     ndi=1.2     UTnbr=207m   lnBr=-23     kbq=85.8u
.PARAM  Wcml={beta4c*4*c}        
.PARAM  aubr={0.93m*UBr}
.PARAM  dvgs={0.1-0.06*Vth0}

.PARAM  f1=80p         f2=54p         f3=204p        f4=320p        f5=390p
.PARAM  U0=0.5         nd=0.42        nc=0.5         g1=4           bb=-1.5
.PARAM  sl=150p        remp=0p        ta=60n         td=20n

.PARAM  Vmin=1.3       Vmax=2.3       dCmax=0.35
.PARAM  Vth={Vth0+(Vmax-Vth0)*limit(dVth,0,1)-(Vmin-Vth0)*limit(dVth,-1,0)}
.PARAM  p0={Wcml*a*((1-f_bet)*(T0/Tref)**mu_bet+f_bet)    }
.PARAM  Rlim={(Rmax-Rs-(Unn-Vth0-Inn*Rs-SQRT((Unn-Vth0-Inn*Rs)**2-4*c*Inn/p0))/(2*c*Inn))/(1+rpa*(Inn/a)**2)} 
.PARAM  dRd={Rd/a+if(dVth==0,limit(dR,0,1)*max(Rlim-Rd/a,0),0)} 
.PARAM  bet={Wcml}

.PARAM  dC1={1+dCmax*limit(dC,0,1)} 
.PARAM  Cox={f1*a*dC1}
.PARAM  Cds0={f2*a*dC1}
.PARAM  Cgs0={f3*a*dC1}
.PARAM  Cox1={f5*a*dC1}
.PARAM  Crand={remp*SQRT(a)}
.PARAM  dRdi={Rdi/a}

.FUNC U1(Uds,T)       {(SQRT(1+4*(0.4+(T-T0-25)*2m)*abs(Uds))-1)/2/(0.4+(T-T0-25)*2m)}
.FUNC I2(p,Uee,z1,pp) {if(Uee>pp,(Uee-c*z1)*z1,p*(pp-p)/c*exp((Uee-pp-(min(0,Uee))**2)/p))}
.FUNC Ig(Uds,T,p,Uee) {bet*((1-f_bet)*(T0/T)**mu_bet+f_bet)*I2(p,Uee,min(Uds,Uee/(2*c)),min(2*p,p+c*Uds))}
.FUNC Iges(Uds,Ugs,T) 
 +{a*(sgn(Uds)*Ig(U1(Uds,T),T,1/(ph0-ph1*T),Ugs-Vth+auth*(T-Tref))+exp(min(lnBr+(abs(Uds)-UBr-aubr*(T-Tref))/UTnbr,25)))}

.FUNC Isjt(Tj)           {exp(min(lnIsj+(Tj/Tref-1)*1.12/(ndi*kbq*Tj),9))*(Tj/Tref)**1.5}
.FUNC Idiode(Usd,Tj,Iss) {exp(min(log(Iss)+Usd/(ndi*kbq*Tj),9))-Iss}
.FUNC Idiod(Usd,Tj)      {a*Idiode(Usd,Tj,Isjt(Tj))}

.FUNC QCdg(x,z)  {if(f4>f5,(f5**2-(f4-z*sl)**2)/(2*sl)+f5*min(x,(f4-f5)/sl),f4*z-sl*z**2/2-f5*max((f4-f5)/sl-x,0))}

E_Edg     d   ox  VALUE {V(d,g)-(min(V(d,g),-bb)+1/(g1*(1-nc))*((1/(1+g1*max(V(d,g)+bb,0)))**(nc-1)-1))}
C_Cdg     ox  g   {Cox}
E_Edg1    d   ox1 VALUE {V(d,g)-QCdg(V(d,g),limit(V(d,g),(f4-f5)/sl,f4/sl))/f5}
C_Cdg1    ox1 g   {Cox1}
C_Cdg2    d   g   {Crand}

E_Eds     d edep  VALUE {(V(d2,s)-I(V_sense3)/Cds0)}
C_Cds  edep    s  {Cds0}
C_Cds2   d2    s  {Cds0/500}

C_Cgs     g    s  {Cgs0}

G_chan    d    s  VALUE={Iges(V(d,s),V(g,s),T0+limit(V(Tj),-200,350))}
E_RMos   d1    d  VALUE={I(V_sense)*(Rf*dRd+(1-Rf)*dRd*((limit(V(Tj),-200,999)+T0)/Tref)**nmu)*(1+rpa*(I(V_sense)/a)**2)}
V_sense  dd   d1  0
G_diode   s   d2  VALUE={Idiod(V(s,d2),T0+limit(V(Tj),-200,499))}
R_Rdio   d2   d3  {dRdi}
V_sense2 d1   d3  0

L_L001    a    c  {td/(ta+td)}
R_R001    a    b  {1/ta}
V_sense3  c    f  0
R_sense3  f    0  1
E_E001    b    0  VALUE {I(V_sense2)}
E_E002    e    0  VALUE {1Meg*Cds0*(1/(1-nd)*U0**nd*(limit(U0+V(d2,s),U0/2,2*UBr))**(1-nd)+2**nd*min(V(d2,s)+U0/2,0))}
R_R002    e    c  1Meg

R1        g    s  1G
Rd01      d    s  500Meg
Rd02     d2    s  500Meg
Rd03     d1    d  10k

G_TH      0    Tj  VALUE = {heat*LIMIT(I(V_sense)*V(dd,s),0,100k)}

.ENDS
*$

**************************************************************************************


.SUBCKT K_600_a_var dd g s Tj PARAMS: a=1 dVth=0 dR=0 dgfs=0 Inn=1 Unn=1 Rmax=1
+gmin=1 Rs=1 Rp=1 dC=0 heat=1

.PARAM  Vth0=2.07      beta4c=0.157   ph0=25.7       ph1=0.038      Ubr=650
.PARAM  Rd=11          nmu=2.7        Rf=0.1         rpa=0.58357    lnIsj=-24.7
.PARAM  Rdi=0.2

.PARAM  Tref=298     T0=273      auth=3m      c=0.82       mu_bet=0.4
.PARAM  f_bet=-2     ndi=1.2     UTnbr=207m   lnBr=-23     kbq=85.8u
.PARAM  Wcml={beta4c*4*c}        
.PARAM  aubr={0.93m*UBr}
.PARAM  dvgs={0.1-0.06*Vth0}

.PARAM  f1=80p         f2=60p         f3=204p        f4=320p        f5=390p
.PARAM  U0=0.5         nd=0.42        nc=0.5         g1=7           bb=-1.5
.PARAM  sl=150p        remp=0p        ta=60n         td=20n

.PARAM  Vmin=1.3       Vmax=2.3       dCmax=0.35
.PARAM  Vth={Vth0+(Vmax-Vth0)*limit(dVth,0,1)-(Vmin-Vth0)*limit(dVth,-1,0)}
.PARAM  p0={Wcml*a*((1-f_bet)*(T0/Tref)**mu_bet+f_bet)    }
.PARAM  Rlim={(Rmax-Rs-(Unn-Vth0-Inn*Rs-SQRT((Unn-Vth0-Inn*Rs)**2-4*c*Inn/p0))/(2*c*Inn))/(1+rpa*(Inn/a)**2)} 
.PARAM  dRd={Rd/a+if(dVth==0,limit(dR,0,1)*max(Rlim-Rd/a,0),0)} 
.PARAM  bet={Wcml}

.PARAM  dC1={1+dCmax*limit(dC,0,1)} 
.PARAM  Cox={f1*a*dC1}
.PARAM  Cds0={f2*a*dC1}
.PARAM  Cgs0={f3*a*dC1}
.PARAM  Cox1={f5*a*dC1}
.PARAM  Crand={remp*SQRT(a)}
.PARAM  dRdi={Rdi/a}

.FUNC U1(Uds,T)       {(SQRT(1+4*(0.4+(T-T0-25)*2m)*abs(Uds))-1)/2/(0.4+(T-T0-25)*2m)}
.FUNC I2(p,Uee,z1,pp) {if(Uee>pp,(Uee-c*z1)*z1,p*(pp-p)/c*exp((Uee-pp-(min(0,Uee))**2)/p))}
.FUNC Ig(Uds,T,p,Uee) {bet*((1-f_bet)*(T0/T)**mu_bet+f_bet)*I2(p,Uee,min(Uds,Uee/(2*c)),min(2*p,p+c*Uds))}
.FUNC Iges(Uds,Ugs,T) 
 +{a*(sgn(Uds)*Ig(U1(Uds,T),T,1/(ph0-ph1*T),Ugs-Vth+auth*(T-Tref))+exp(min(lnBr+(abs(Uds)-UBr-aubr*(T-Tref))/UTnbr,25)))}

.FUNC Isjt(Tj)           {exp(min(lnIsj+(Tj/Tref-1)*1.12/(ndi*kbq*Tj),9))*(Tj/Tref)**1.5}
.FUNC Idiode(Usd,Tj,Iss) {exp(min(log(Iss)+Usd/(ndi*kbq*Tj),9))-Iss}
.FUNC Idiod(Usd,Tj)      {a*Idiode(Usd,Tj,Isjt(Tj))}

.FUNC QCdg(x,z)  {if(f4>f5,(f5**2-(f4-z*sl)**2)/(2*sl)+f5*min(x,(f4-f5)/sl),f4*z-sl*z**2/2-f5*max((f4-f5)/sl-x,0))}

E_Edg     d   ox  VALUE {V(d,g)-(min(V(d,g),-bb)+1/(g1*(1-nc))*((1/(1+g1*max(V(d,g)+bb,0)))**(nc-1)-1))}
C_Cdg     ox  g   {Cox}
E_Edg1    d   ox1 VALUE {V(d,g)-QCdg(V(d,g),limit(V(d,g),(f4-f5)/sl,f4/sl))/f5}
C_Cdg1    ox1 g   {Cox1}
C_Cdg2    d   g   {Crand}

E_Eds     d edep  VALUE {(V(d2,s)-I(V_sense3)/Cds0)}
C_Cds  edep    s  {Cds0}
C_Cds2   d2    s  {Cds0/500}

C_Cgs     g    s  {Cgs0}

G_chan    d    s  VALUE={Iges(V(d,s),V(g,s),T0+limit(V(Tj),-200,350))}
E_RMos   d1    d  VALUE={I(V_sense)*(Rf*dRd+(1-Rf)*dRd*((limit(V(Tj),-200,999)+T0)/Tref)**nmu)*(1+rpa*(I(V_sense)/a)**2)}
V_sense  dd   d1  0
G_diode   s   d2  VALUE={Idiod(V(s,d2),T0+limit(V(Tj),-200,499))}
R_Rdio   d2   d3  {dRdi}
V_sense2 d1   d3  0

L_L001    a    c  {td/(ta+td)}
R_R001    a    b  {1/ta}
V_sense3  c    f  0
R_sense3  f    0  1
E_E001    b    0  VALUE {I(V_sense2)}
E_E002    e    0  VALUE {1Meg*Cds0*(1/(1-nd)*U0**nd*(limit(U0+V(d2,s),U0/2,2*UBr))**(1-nd)+2**nd*min(V(d2,s)+U0/2,0))}
R_R002    e    c  1Meg

R1        g    s  1G
Rd01      d    s  500Meg
Rd02     d2    s  500Meg
Rd03     d1    d  20k

G_TH      0    Tj  VALUE = {heat*LIMIT(I(V_sense)*V(dd,s),0,100k)}

.ENDS
*$

**************************************************************************************


.SUBCKT K_600_d_var dd g s Tj PARAMS: a=1 dVth=0 dR=0 dgfs=0 Inn=1 Unn=1 Rmax=1
+gmin=1 Rs=1 Rp=1 dC=0 heat=1

.PARAM  Vth0=-1.15     beta4c=0.157   ph0=20         ph1=0.026      Ubr=650
.PARAM  Rd=11          nmu=2.7        Rf=0.1         rpa=0.58357    lnIsj=-24.7
.PARAM  Rdi=0.2

.PARAM  Tref=298     T0=273      auth=3m      c=0.82       mu_bet=0.4
.PARAM  f_bet=-2     ndi=1.2     UTnbr=207m   lnBr=-23     kbq=85.8u
.PARAM  Wcml={beta4c*4*c}        
.PARAM  aubr={0.93m*UBr}
.PARAM  dvgs={0.1-0.06*Vth0}

.PARAM  f1=100p        f2=60p         f3=204p        f4=435p        f5=355p
.PARAM  U0=0.5         nd=0.43        nc=0.5         g1=9           bb=-9.8
.PARAM  sl=37p         remp=0p        ta=100n        td=30n

.PARAM  Vmin=-2.1      Vmax=-1        dCmax=0.35
.PARAM  Vth={Vth0+(Vmax-Vth0)*limit(dVth,0,1)-(Vmin-Vth0)*limit(dVth,-1,0)}
.PARAM  p0={Wcml*a*((1-f_bet)*(T0/Tref)**mu_bet+f_bet)    }
.PARAM  Rlim={(Rmax-Rs-(Unn-Vth0-Inn*Rs-SQRT((Unn-Vth0-Inn*Rs)**2-4*c*Inn/p0))/(2*c*Inn))/(1+rpa*(Inn/a)**2)} 
.PARAM  dRd={Rd/a+if(dVth==0,limit(dR,0,1)*max(Rlim-Rd/a,0),0)} 
.PARAM  bet={Wcml}

.PARAM  dC1={1+dCmax*limit(dC,0,1)} 
.PARAM  Cox={f1*a*dC1}
.PARAM  Cds0={f2*a*dC1}
.PARAM  Cgs0={f3*a*dC1}
.PARAM  Cox1={f5*a*dC1}
.PARAM  Crand={remp*SQRT(a)}
.PARAM  dRdi={Rdi/a}

.FUNC U1(Uds,T)       {(SQRT(1+4*(0.4+(T-T0-25)*2m)*abs(Uds))-1)/2/(0.4+(T-T0-25)*2m)}
.FUNC I2(p,Uee,z1,pp) {if(Uee>pp,(Uee-c*z1)*z1,p*(pp-p)/c*exp((Uee-pp-(min(0,Uee))**2)/p))}
.FUNC Ig(Uds,T,p,Uee) {bet*((1-f_bet)*(T0/T)**mu_bet+f_bet)*I2(p,Uee,min(Uds,Uee/(2*c)),min(2*p,p+c*Uds))}
.FUNC Iges(Uds,Ugs,T) 
 +{a*(sgn(Uds)*Ig(U1(Uds,T),T,1/(ph0-ph1*T),Ugs-Vth+auth*(T-Tref))+exp(min(lnBr+(abs(Uds)-UBr-aubr*(T-Tref))/UTnbr,25)))}

.FUNC Isjt(Tj)           {exp(min(lnIsj+(Tj/Tref-1)*1.12/(ndi*kbq*Tj),9))*(Tj/Tref)**1.5}
.FUNC Idiode(Usd,Tj,Iss) {exp(min(log(Iss)+Usd/(ndi*kbq*Tj),9))-Iss}
.FUNC Idiod(Usd,Tj)      {a*Idiode(Usd,Tj,Isjt(Tj))}

.FUNC QCdg(x,z)  {if(f4>f5,(f5**2-(f4-z*sl)**2)/(2*sl)+f5*min(x,(f4-f5)/sl),f4*z-sl*z**2/2-f5*max((f4-f5)/sl-x,0))}

E_Edg     d   ox  VALUE {V(d,g)-(min(V(d,g),-bb)+1/(g1*(1-nc))*((1/(1+g1*max(V(d,g)+bb,0)))**(nc-1)-1))}
C_Cdg     ox  g   {Cox}
E_Edg1    d   ox1 VALUE {V(d,g)-QCdg(V(d,g),limit(V(d,g),(f4-f5)/sl,f4/sl))/f5}
C_Cdg1    ox1 g   {Cox1}
C_Cdg2    d   g   {Crand}

E_Eds     d edep  VALUE {(V(d2,s)-I(V_sense3)/Cds0)}
C_Cds  edep    s  {Cds0}
C_Cds2   d2    s  {Cds0/500}

C_Cgs     g    s  {Cgs0}

G_chan    d    s  VALUE={Iges(V(d,s),V(g,s),T0+limit(V(Tj),-200,350))}
E_RMos   d1    d  VALUE={I(V_sense)*(Rf*dRd+(1-Rf)*dRd*((limit(V(Tj),-200,999)+T0)/Tref)**nmu)*(1+rpa*(I(V_sense)/a)**2)}
V_sense  dd   d1  0
G_diode   s   d2  VALUE={Idiod(V(s,d2),T0+limit(V(Tj),-200,499))}
R_Rdio   d2   d3  {dRdi}
V_sense2 d1   d3  0

L_L001    a    c  {td/(ta+td)}
R_R001    a    b  {1/ta}
V_sense3  c    f  0
R_sense3  f    0  1
E_E001    b    0  VALUE {I(V_sense2)}
E_E002    e    0  VALUE {1Meg*Cds0*(1/(1-nd)*U0**nd*(limit(U0+V(d2,s),U0/2,2*UBr))**(1-nd)+2**nd*min(V(d2,s)+U0/2,0))}
R_R002    e    c  1Meg

R1        g    s  1G
Rd01      d    s  500Meg
Rd02     d2    s  500Meg
Rd03     d1    d  20k

G_TH      0    Tj  VALUE = {heat*LIMIT(I(V_sense)*V(dd,s),0,100k)}

.ENDS
*$

**************************************************************************************


.SUBCKT K_600_e_var dd g s Tj PARAMS: a=1 dVth=0 dR=0 dgfs=0 Inn=1 Unn=1 Rmax=1
+gmin=1 Rs=1 Rp=1 dC=0 heat=1

.PARAM  Vth0=-1.75     beta4c=0.206   ph0=20         ph1=0.026      Ubr=650
.PARAM  Rd=11          nmu=2.7        Rf=0.1         rpa=0.58357    lnIsj=-24.7
.PARAM  Rdi=0.2

.PARAM  Tref=298     T0=273      auth=3m      c=0.82       mu_bet=0.4
.PARAM  f_bet=-2     ndi=1.2     UTnbr=207m   lnBr=-23     kbq=85.8u
.PARAM  Wcml={beta4c*4*c}        
.PARAM  aubr={0.93m*UBr}
.PARAM  dvgs={0.1-0.06*Vth0}

.PARAM  f1=100p        f2=100p        f3=500p        f4=435p        f5=500p
.PARAM  U0=0.5         nd=0.4         nc=0.5         g1=9           bb=-9.8
.PARAM  sl=37p         remp=2p        ta=60n         td=20n

.PARAM  Vmin=-2.7      Vmax=-1.6      dCmax=0.35
.PARAM  Vth={Vth0+(Vmax-Vth0)*limit(dVth,0,1)-(Vmin-Vth0)*limit(dVth,-1,0)}
.PARAM  p0={Wcml*a*((1-f_bet)*(T0/Tref)**mu_bet+f_bet)    }
.PARAM  Rlim={(Rmax-Rs-(Unn-Vth0-Inn*Rs-SQRT((Unn-Vth0-Inn*Rs)**2-4*c*Inn/p0))/(2*c*Inn))/(1+rpa*(Inn/a)**2)} 
.PARAM  dRd={Rd/a+if(dVth==0,limit(dR,0,1)*max(Rlim-Rd/a,0),0)} 
.PARAM  bet={Wcml}

.PARAM  dC1={1+dCmax*limit(dC,0,1)} 
.PARAM  Cox={f1*a*dC1}
.PARAM  Cds0={f2*a*dC1}
.PARAM  Cgs0={f3*a*dC1}
.PARAM  Cox1={f5*a*dC1}
.PARAM  Crand={remp*SQRT(a)}
.PARAM  dRdi={Rdi/a}

.FUNC U1(Uds,T)       {(SQRT(1+4*(0.4+(T-T0-25)*2m)*abs(Uds))-1)/2/(0.4+(T-T0-25)*2m)}
.FUNC I2(p,Uee,z1,pp) {if(Uee>pp,(Uee-c*z1)*z1,p*(pp-p)/c*exp((Uee-pp-(min(0,Uee))**2)/p))}
.FUNC Ig(Uds,T,p,Uee) {bet*((1-f_bet)*(T0/T)**mu_bet+f_bet)*I2(p,Uee,min(Uds,Uee/(2*c)),min(2*p,p+c*Uds))}
.FUNC Iges(Uds,Ugs,T) 
 +{a*(sgn(Uds)*Ig(U1(Uds,T),T,1/(ph0-ph1*T),Ugs-Vth+auth*(T-Tref))+exp(min(lnBr+(abs(Uds)-UBr-aubr*(T-Tref))/UTnbr,25)))}

.FUNC Isjt(Tj)           {exp(min(lnIsj+(Tj/Tref-1)*1.12/(ndi*kbq*Tj),9))*(Tj/Tref)**1.5}
.FUNC Idiode(Usd,Tj,Iss) {exp(min(log(Iss)+Usd/(ndi*kbq*Tj),9))-Iss}
.FUNC Idiod(Usd,Tj)      {a*Idiode(Usd,Tj,Isjt(Tj))}

.FUNC QCdg(x,z)  {if(f4>f5,(f5**2-(f4-z*sl)**2)/(2*sl)+f5*min(x,(f4-f5)/sl),f4*z-sl*z**2/2-f5*max((f4-f5)/sl-x,0))}

E_Edg     d   ox  VALUE {V(d,g)-(min(V(d,g),-bb)+1/(g1*(1-nc))*((1/(1+g1*max(V(d,g)+bb,0)))**(nc-1)-1))}
C_Cdg     ox  g   {Cox}
E_Edg1    d   ox1 VALUE {V(d,g)-QCdg(V(d,g),limit(V(d,g),(f4-f5)/sl,f4/sl))/f5}
C_Cdg1    ox1 g   {Cox1}
C_Cdg2    d   g   {Crand}

E_Eds     d edep  VALUE {(V(d2,s)-I(V_sense3)/Cds0)}
C_Cds  edep    s  {Cds0}
C_Cds2   d2    s  {Cds0/500}

C_Cgs     g    s  {Cgs0}

G_chan    d    s  VALUE={Iges(V(d,s),V(g,s),T0+limit(V(Tj),-200,350))}
E_RMos   d1    d  VALUE={I(V_sense)*(Rf*dRd+(1-Rf)*dRd*((limit(V(Tj),-200,999)+T0)/Tref)**nmu)*(1+rpa*(I(V_sense)/a)**2)}
V_sense  dd   d1  0
G_diode   s   d2  VALUE={Idiod(V(s,d2),T0+limit(V(Tj),-200,499))}
R_Rdio   d2   d3  {dRdi}
V_sense2 d1   d3  0

L_L001    a    c  {td/(ta+td)}
R_R001    a    b  {1/ta}
V_sense3  c    f  0
R_sense3  f    0  1
E_E001    b    0  VALUE {I(V_sense2)}
E_E002    e    0  VALUE {1Meg*Cds0*(1/(1-nd)*U0**nd*(limit(U0+V(d2,s),U0/2,2*UBr))**(1-nd)+2**nd*min(V(d2,s)+U0/2,0))}
R_R002    e    c  1Meg

R1        g    s  1G
Rd01      d    s  500Meg
Rd02     d2    s  500Meg
Rd03     d1    d  100k

G_TH      0    Tj  VALUE = {heat*LIMIT(I(V_sense)*V(dd,s),0,100k)}

.ENDS
*$



.SUBCKT BSS131 drain gate source Tj Tcase PARAMS: dVth=0 dRdson=0 dgfs=0 dC=0 Zthtype=0

.PARAM Rs=0.074     Rg=10        Ls=3n        Ld=1n        Lg=3n
.PARAM Inn=0.1      Unn=10       Rmax=14
.PARAM act=0.28

X1  d1 g s Tj K_240_a_var PARAMS: a={act} dVth={dVth} dR={dRdson} Inn={Inn} Unn={Unn} 
                                        +Rmax={Rmax} dgfs={dgfs} Rs={Rs} dC={dC} heat=1

Rg    g1     g    {Rg}   
Lg    gate   g1   {Lg*if(dgfs==99,0,1)}
Gs    s1     s    VALUE={V(s1,s)/(Rs*(1+(limit(V(Tj),-200,999)-25)*4m))}
Rsa   s1     s    1Meg
Ls    source s1   {Ls*if(dgfs==99,0,1)}
Ld    drain  d1   {Ld*if(dgfs==99,0,1)}

Rth1  Tj      t1              {624.77m+limit(Zthtype,0,1)*231.23m}
Rth2  t1      t2              {2.85+limit(Zthtype,0,1)*1.06}
Rth3  t2      t3              {5.96+limit(Zthtype,0,1)*781.17m}
Rth4  t3      t4              {68.15+limit(Zthtype,0,1)*58.03}
Rth5  t4      Tcase           {79.56+limit(Zthtype,0,1)*67.75}
Cth1  Tj      0               10.376u
Cth2  t1      0               17.965u
Cth3  t2      0               180.456u
Cth4  t3      0               374.154u
Cth5  t4      0               4.696m


.ENDS
*$

********************

.SUBCKT BSS87 drain gate source Tj Tcase PARAMS: dVth=0 dRdson=0 dgfs=0 dC=0 Zthtype=0

.PARAM Rs=0.082     Rg=10        Ls=3n        Ld=1n        Lg=3n
.PARAM Inn=0.26     Unn=10       Rmax=6
.PARAM act=0.54

X1  d1 g s Tj K_240_b_var PARAMS: a={act} dVth={dVth} dR={dRdson} Inn={Inn} Unn={Unn} 
                                        +Rmax={Rmax} dgfs={dgfs} Rs={Rs} dC={dC} heat=1

Rg    g1     g    {Rg}   
Lg    gate   g1   {Lg*if(dgfs==99,0,1)}
Gs    s1     s    VALUE={V(s1,s)/(Rs*(1+(limit(V(Tj),-200,999)-25)*4m))}
Rsa   s1     s    1Meg
Ls    source s1   {Ls*if(dgfs==99,0,1)}
Ld    drain  d1   {Ld*if(dgfs==99,0,1)}

Rth1  Tj      t1              {166.55m+limit(Zthtype,0,1)*61.64m}
Rth2  t1      t2              {730.55m+limit(Zthtype,0,1)*270.37m}
Rth3  t2      t3              {2.71+limit(Zthtype,0,1)*733.69m}
Rth4  t3      t4              {605m+limit(Zthtype,0,1)*2.11}
Rth5  t4      Tcase           {581m+limit(Zthtype,0,1)*2.03}
Cth1  Tj      0               13.4u
Cth2  t1      0               7.5u
Cth3  t2      0               43.4u
Cth4  t3      0               400u
Cth5  t4      0               600u
Cth6  Tcase   0               4m

.ENDS
*$

********************

.SUBCKT BSP89 drain gate source Tj Tcase PARAMS: dVth=0 dRdson=0 dgfs=0 dC=0 Zthtype=0

.PARAM Rs=0.027     Rg=10        Ls=3n        Ld=1n        Lg=3n
.PARAM Inn=0.35     Unn=10       Rmax=6
.PARAM act=0.54

X1  d1 g s Tj K_240_b_var PARAMS: a={act} dVth={dVth} dR={dRdson} Inn={Inn} Unn={Unn} 
                                        +Rmax={Rmax} dgfs={dgfs} Rs={Rs} dC={dC} heat=1

Rg    g1     g    {Rg}   
Lg    gate   g1   {Lg*if(dgfs==99,0,1)}
Gs    s1     s    VALUE={V(s1,s)/(Rs*(1+(limit(V(Tj),-200,999)-25)*4m))}
Rsa   s1     s    1Meg
Ls    source s1   {Ls*if(dgfs==99,0,1)}
Ld    drain  d1   {Ld*if(dgfs==99,0,1)}

Rth1  Tj      t1              {166.55m+limit(Zthtype,0,1)*61.64m}
Rth2  t1      t2              {730.55m+limit(Zthtype,0,1)*270.37m}
Rth3  t2      t3              {7.81+limit(Zthtype,0,1)*741.69m}
Rth4  t3      t4              {7.4+limit(Zthtype,0,1)*9.35m}
Rth5  t4      Tcase           {7.8+limit(Zthtype,0,1)*9.85m}
Cth1  Tj      0               13.4u
Cth2  t1      0               7.5u
Cth3  t2      0               149.668u
Cth4  t3      0               1.95m
Cth5  t4      0               48.845m


.ENDS
*$

********************

.SUBCKT BSP88 drain gate source Tj Tcase PARAMS: dVth=0 dRdson=0 dgfs=0 dC=0 Zthtype=0

.PARAM Rs=0.027     Rg=10        Ls=3n        Ld=1n        Lg=3n
.PARAM Inn=0.35     Unn=10       Rmax=6
.PARAM act=0.54

X1  d1 g s Tj K_240_c_var PARAMS: a={act} dVth={dVth} dR={dRdson} Inn={Inn} Unn={Unn} 
                                        +Rmax={Rmax} dgfs={dgfs} Rs={Rs} dC={dC} heat=1

Rg    g1     g    {Rg}   
Lg    gate   g1   {Lg*if(dgfs==99,0,1)}
Gs    s1     s    VALUE={V(s1,s)/(Rs*(1+(limit(V(Tj),-200,999)-25)*4m))}
Rsa   s1     s    1Meg
Ls    source s1   {Ls*if(dgfs==99,0,1)}
Ld    drain  d1   {Ld*if(dgfs==99,0,1)}

Rth1  Tj      t1              {166.55m+limit(Zthtype,0,1)*61.64m}
Rth2  t1      t2              {730.55m+limit(Zthtype,0,1)*270.37m}
Rth3  t2      t3              {7.81+limit(Zthtype,0,1)*741.69m}
Rth4  t3      t4              {7.4+limit(Zthtype,0,1)*9.35m}
Rth5  t4      Tcase           {7.8+limit(Zthtype,0,1)*9.85m}
Cth1  Tj      0               13.4u
Cth2  t1      0               7.5u
Cth3  t2      0               149.668u
Cth4  t3      0               1.95m
Cth5  t4      0               48.845m


.ENDS
*$

********************

.SUBCKT BSP129 drain gate source Tj Tcase PARAMS: dVth=0 dRdson=0 dgfs=0 dC=0 Zthtype=0

.PARAM Rs=0.027     Rg=10        Ls=3n        Ld=1n        Lg=3n
.PARAM Inn=0.025    Unn=0        Rmax=20
.PARAM act=0.54

X1  d1 g s Tj K_240_d_var PARAMS: a={act} dVth={dVth} dR={dRdson} Inn={Inn} Unn={Unn} 
                                        +Rmax={Rmax} dgfs={dgfs} Rs={Rs} dC={dC} heat=1

Rg    g1     g    {Rg}   
Lg    gate   g1   {Lg*if(dgfs==99,0,1)}
Gs    s1     s    VALUE={V(s1,s)/(Rs*(1+(limit(V(Tj),-200,999)-25)*4m))}
Rsa   s1     s    1Meg
Ls    source s1   {Ls*if(dgfs==99,0,1)}
Ld    drain  d1   {Ld*if(dgfs==99,0,1)}

Rth1  Tj      t1              {166.55m+limit(Zthtype,0,1)*61.64m}
Rth2  t1      t2              {730.55m+limit(Zthtype,0,1)*270.37m}
Rth3  t2      t3              {7.81+limit(Zthtype,0,1)*741.69m}
Rth4  t3      t4              {7.4+limit(Zthtype,0,1)*9.35m}
Rth5  t4      Tcase           {7.8+limit(Zthtype,0,1)*9.85m}
Cth1  Tj      0               13.4u
Cth2  t1      0               7.5u
Cth3  t2      0               149.668u
Cth4  t3      0               1.95m
Cth5  t4      0               48.845m


.ENDS
*$

********************

.SUBCKT SISC0_97N24D drain gate source Tj Tcase PARAMS: dVth=0 dRdson=0 dgfs=0 dC=0 Zthtype=0

.PARAM Rs=0.005     Rg=10      
.PARAM Inn=0.025    Unn=0        Rmax=20
.PARAM act=0.54

X1  drain g s Tj K_240_d_var PARAMS: a={act} dVth={dVth} dR={dRdson} Inn={Inn} Unn={Unn} 
                                        +Rmax={Rmax} dgfs={dgfs} Rs={Rs} dC={dC} heat=1

Rg    gate     g    {Rg}   

Gs    source     s    VALUE={V(source,s)/(Rs*(1+(limit(V(Tj),-200,999)-25)*4m))}
Rsa   source     s    1Meg



Rth1  Tj      t1              {166.55m+limit(Zthtype,0,1)*61.64m}
Rth2  t1      t2              {730.55m+limit(Zthtype,0,1)*270.37m}
Rth3  t2      t3              {2+limit(Zthtype,0,1)*741.69m}
Rth4  t3      t4              {1p+limit(Zthtype,0,1)*0p}
Rth5  t4      Tcase           {1p+limit(Zthtype,0,1)*0p}
Cth1  Tj      0               13.4u
Cth2  t1      0               7.5u
Cth3  t2      0               149.668u
Cth4  t3      0               1p
Cth5  t4      0               1p


.ENDS

********************

.SUBCKT BSS139 drain gate source Tj Tcase PARAMS: dVth=0 dRdson=0 dgfs=0 dC=0 Zthtype=0

.PARAM Rs=0.074     Rg=10        Ls=3n        Ld=1n        Lg=3n
.PARAM Inn=0.015    Unn=0        Rmax=30
.PARAM act=0.28

X1  d1 g s Tj K_250_d_var PARAMS: a={act} dVth={dVth} dR={dRdson} Inn={Inn} Unn={Unn} 
                                        +Rmax={Rmax} dgfs={dgfs} Rs={Rs} dC={dC} heat=1

Rg    g1     g    {Rg}   
Lg    gate   g1   {Lg*if(dgfs==99,0,1)}
Gs    s1     s    VALUE={V(s1,s)/(Rs*(1+(limit(V(Tj),-200,999)-25)*4m))}
Rsa   s1     s    1Meg
Ls    source s1   {Ls*if(dgfs==99,0,1)}
Ld    drain  d1   {Ld*if(dgfs==99,0,1)}

Rth1  Tj      t1              {624.77m+limit(Zthtype,0,1)*231.23m}
Rth2  t1      t2              {2.85+limit(Zthtype,0,1)*1.06}
Rth3  t2      t3              {5.96+limit(Zthtype,0,1)*781.17m}
Rth4  t3      t4              {68.15+limit(Zthtype,0,1)*58.03}
Rth5  t4      Tcase           {79.56+limit(Zthtype,0,1)*67.75}
Cth1  Tj      0               10.376u
Cth2  t1      0               17.965u
Cth3  t2      0               180.456u
Cth4  t3      0               374.154u
Cth5  t4      0               4.696m


.ENDS
*$

********************

.SUBCKT BSP324 drain gate source Tj Tcase PARAMS: dVth=0 dRdson=0 dgfs=0 dC=0 Zthtype=0

.PARAM Rs=0.027     Rg=10        Ls=3n        Ld=1n        Lg=3n
.PARAM Inn=0.17     Unn=10       Rmax=25
.PARAM act=0.47

X1  d1 g s Tj K_400_a_var PARAMS: a={act} dVth={dVth} dR={dRdson} Inn={Inn} Unn={Unn} 
                                        +Rmax={Rmax} dgfs={dgfs} Rs={Rs} dC={dC} heat=1

Rg    g1     g    {Rg}   
Lg    gate   g1   {Lg*if(dgfs==99,0,1)}
Gs    s1     s    VALUE={V(s1,s)/(Rs*(1+(limit(V(Tj),-200,999)-25)*4m))}
Rsa   s1     s    1Meg
Ls    source s1   {Ls*if(dgfs==99,0,1)}
Ld    drain  d1   {Ld*if(dgfs==99,0,1)}

Rth1  Tj      t1              {685.56m+limit(Zthtype,0,1)*253.73m}
Rth2  t1      t2              {2.03+limit(Zthtype,0,1)*756.67m}
Rth3  t2      t3              {5.71+limit(Zthtype,0,1)*221.88m}
Rth4  t3      t4              {5.53+limit(Zthtype,0,1)*810.97m}
Rth5  t4      Tcase           {7.85+limit(Zthtype,0,1)*1.15}
Cth1  Tj      0               23.846u
Cth2  t1      0               48.38u
Cth3  t2      0               177.844u
Cth4  t3      0               1.642m
Cth5  t4      0               48.845m


.ENDS
*$

********************

.SUBCKT SISC1_4N40E drain gate source Tj Tcase PARAMS: dVth=0 dRdson=0 dgfs=0 dC=0 Zthtype=0

.PARAM Rs=0.005     Rg=10        
.PARAM Inn=0.17     Unn=10       Rmax=25
.PARAM act=0.47

X1  drain g s Tj K_400_a_var PARAMS: a={act} dVth={dVth} dR={dRdson} Inn={Inn} Unn={Unn} 
                                        +Rmax={Rmax} dgfs={dgfs} Rs={Rs} dC={dC} heat=1

Rg    gate     g    {Rg}   

Gs    source     s    VALUE={V(source,s)/(Rs*(1+(limit(V(Tj),-200,999)-25)*4m))}
Rsa   source     s    1Meg



Rth1  Tj      t1              {685.56m+limit(Zthtype,0,1)*253.73m}
Rth2  t1      t2              {2.03+limit(Zthtype,0,1)*756.67m}
Rth3  t2      t3              {624.96m+limit(Zthtype,0,1)*222.92m}
Rth4  t3      t4              {1p+limit(Zthtype,0,1)*0}
Rth5  t4      Tcase           {1p+limit(Zthtype,0,1)*0}
Cth1  Tj      0               23.846u
Cth2  t1      0               48.38u
Cth3  t2      0               177.844u
Cth4  t3      0               1p
Cth5  t4      0               1p


.ENDS
*$

********************

.SUBCKT BSP125 drain gate source Tj Tcase PARAMS: dVth=0 dRdson=0 dgfs=0 dC=0 Zthtype=0

.PARAM Rs=0.027     Rg=10        Ls=3n        Ld=1n        Lg=3n
.PARAM Inn=0.12     Unn=10       Rmax=45
.PARAM act=0.47

X1  d1 g s Tj K_600_a_var PARAMS: a={act} dVth={dVth} dR={dRdson} Inn={Inn} Unn={Unn} 
                                        +Rmax={Rmax} dgfs={dgfs} Rs={Rs} dC={dC} heat=1

Rg    g1     g    {Rg}   
Lg    gate   g1   {Lg*if(dgfs==99,0,1)}
Gs    s1     s    VALUE={V(s1,s)/(Rs*(1+(limit(V(Tj),-200,999)-25)*4m))}
Rsa   s1     s    1Meg
Ls    source s1   {Ls*if(dgfs==99,0,1)}
Ld    drain  d1   {Ld*if(dgfs==99,0,1)}

Rth1  Tj      t1              {685.56m+limit(Zthtype,0,1)*253.73m}
Rth2  t1      t2              {2.03+limit(Zthtype,0,1)*756.67m}
Rth3  t2      t3              {5.71+limit(Zthtype,0,1)*221.88m}
Rth4  t3      t4              {5.53+limit(Zthtype,0,1)*810.97m}
Rth5  t4      Tcase           {7.85+limit(Zthtype,0,1)*1.15}
Cth1  Tj      0               23.846u
Cth2  t1      0               48.38u
Cth3  t2      0               177.844u
Cth4  t3      0               1p
Cth5  t4      0               1p


.ENDS
*$

********************

.SUBCKT BSS225 drain gate source Tj Tcase PARAMS: dVth=0 dRdson=0 dgfs=0 dC=0 Zthtype=0

.PARAM Rs=0.027     Rg=10        Ls=3n        Ld=1n        Lg=3n
.PARAM Inn=0.12     Unn=10       Rmax=45
.PARAM act=0.47

X1  d1 g s Tj K_600_a_var PARAMS: a={act} dVth={dVth} dR={dRdson} Inn={Inn} Unn={Unn} 
                                        +Rmax={Rmax} dgfs={dgfs} Rs={Rs} dC={dC} heat=1

Rg    g1     g    {Rg}   
Lg    gate   g1   {Lg*if(dgfs==99,0,1)}
Gs    s1     s    VALUE={V(s1,s)/(Rs*(1+(limit(V(Tj),-200,999)-25)*4m))}
Rsa   s1     s    1Meg
Ls    source s1   {Ls*if(dgfs==99,0,1)}
Ld    drain  d1   {Ld*if(dgfs==99,0,1)}

Rth1  Tj      t1              {166.55m+limit(Zthtype,0,1)*61.64m}
Rth2  t1      t2              {730.55m+limit(Zthtype,0,1)*270.37m}
Rth3  t2      t3              {2.8+limit(Zthtype,0,1)*892.38m}
Rth4  t3      t4              {605m+limit(Zthtype,0,1)*1.99}
Rth5  t4      Tcase           {581m+limit(Zthtype,0,1)*1.91}
Cth1  Tj      0               13.4u
Cth2  t1      0               7.5u
Cth3  t2      0               43.4u
Cth4  t3      0               400u
Cth5  t4      0               600u
Cth6  Tcase   0               4m

.ENDS

********************

.SUBCKT BSS127 drain gate source Tj Tcase PARAMS: dVth=0 dRdson=0 dgfs=0 dC=0 Zthtype=0

.PARAM Rs=0.074     Rg=10        Ls=3n        Ld=1n        Lg=3n
.PARAM Inn=0.016    Unn=10       Rmax=500
.PARAM act=0.04

X1  d1 g s Tj K_600_a_var PARAMS: a={act} dVth={dVth} dR={dRdson} Inn={Inn} Unn={Unn} 
                                        +Rmax={Rmax} dgfs={dgfs} Rs={Rs} dC={dC} heat=1

Rg    g1     g    {Rg}   
Lg    gate   g1   {Lg*if(dgfs==99,0,1)}
Gs    s1     s    VALUE={V(s1,s)/(Rs*(1+(limit(V(Tj),-200,999)-25)*4m))}
Rsa   s1     s    1Meg
Ls    source s1   {Ls*if(dgfs==99,0,1)}
Ld    drain  d1   {Ld*if(dgfs==99,0,1)}

Rth1  Tj      t1              {1.05+limit(Zthtype,0,1)*384.82m}
Rth2  t1      t2              {2.97+limit(Zthtype,0,1)*1.09}
Rth3  t2      t3              {14.08+limit(Zthtype,0,1)*12.96}
Rth4  t3      t4              {47.48+limit(Zthtype,0,1)*18.38}
Rth5  t4      Tcase           {30+limit(Zthtype,0,1)*11.61}
Cth1  Tj      0               3.5u
Cth2  t1      0               1.04u
Cth3  t2      0               1.95u
Cth4  t3      0               414u
Cth5  t4      0               6.75m


.ENDS

********************

.SUBCKT BSP135 drain gate source Tj Tcase PARAMS: dVth=0 dRdson=0 dgfs=0 dC=0 Zthtype=0

.PARAM Rs=0.027     Rg=10        Ls=3n        Ld=1n        Lg=3n
.PARAM Inn=0.01     Unn=0        Rmax=60
.PARAM act=0.47

X1  d1 g s Tj K_600_d_var PARAMS: a={act} dVth={dVth} dR={dRdson} Inn={Inn} Unn={Unn} 
                                        +Rmax={Rmax} dgfs={dgfs} Rs={Rs} dC={dC} heat=1

Rg    g1     g    {Rg}   
Lg    gate   g1   {Lg*if(dgfs==99,0,1)}
Gs    s1     s    VALUE={V(s1,s)/(Rs*(1+(limit(V(Tj),-200,999)-25)*4m))}
Rsa   s1     s    1Meg
Ls    source s1   {Ls*if(dgfs==99,0,1)}
Ld    drain  d1   {Ld*if(dgfs==99,0,1)}

Rth1  Tj      t1              {685.56m+limit(Zthtype,0,1)*253.73m}
Rth2  t1      t2              {2.03+limit(Zthtype,0,1)*756.67m}
Rth3  t2      t3              {5.71+limit(Zthtype,0,1)*221.88m}
Rth4  t3      t4              {5.53+limit(Zthtype,0,1)*810.97m}
Rth5  t4      Tcase           {7.85+limit(Zthtype,0,1)*1.15}
Cth1  Tj      0               44.039u
Cth2  t1      0               43.949u
Cth3  t2      0               360.599u
Cth4  t3      0               6.76m
Cth5  t4      0               103.014m


.ENDS
*$

********************

.SUBCKT SISC1_4N60D drain gate source Tj Tcase PARAMS: dVth=0 dRdson=0 dgfs=0 dC=0 Zthtype=0

.PARAM Rs=0.005     Rg=10        
.PARAM Inn=0.01     Unn=0        Rmax=60
.PARAM act=0.47

X1  drain g s Tj K_600_d_var PARAMS: a={act} dVth={dVth} dR={dRdson} Inn={Inn} Unn={Unn} 
                                        +Rmax={Rmax} dgfs={dgfs} Rs={Rs} dC={dC} heat=1

Rg    gate     g    {Rg}   

Gs    source     s    VALUE={V(source,s)/(Rs*(1+(limit(V(Tj),-200,999)-25)*4m))}
Rsa   source     s    1Meg



Rth1  Tj      t1              {685.56m+limit(Zthtype,0,1)*253.73m}
Rth2  t1      t2              {2.03+limit(Zthtype,0,1)*756.67m}
Rth3  t2      t3              {624.96m+limit(Zthtype,0,1)*222.92m}
Rth4  t3      t4              {1p+limit(Zthtype,0,1)*0}
Rth5  t4      Tcase           {1p+limit(Zthtype,0,1)*0}
Cth1  Tj      0               23.846u
Cth2  t1      0               48.38u
Cth3  t2      0               177.844u
Cth4  t3      0               1p
Cth5  t4      0               1p


.ENDS
*$

********************

.SUBCKT BSS126 drain gate source Tj Tcase PARAMS: dVth=0 dRdson=0 dgfs=0 dC=0 Zthtype=0

.PARAM Rs=0.074     Rg=0.9       Ls=3n        Ld=1n        Lg=3n
.PARAM Inn=0.003    Unn=0        Rmax=700
.PARAM act=0.04

X1  d1 g s Tj K_600_e_var PARAMS: a={act} dVth={dVth} dR={dRdson} Inn={Inn} Unn={Unn} 
                                        +Rmax={Rmax} dgfs={dgfs} Rs={Rs} dC={dC} heat=1

Rg    g1     g    {Rg}   
Lg    gate   g1   {Lg*if(dgfs==99,0,1)}
Gs    s1     s    VALUE={V(s1,s)/(Rs*(1+(limit(V(Tj),-200,999)-25)*4m))}
Rsa   s1     s    1Meg
Ls    source s1   {Ls*if(dgfs==99,0,1)}
Ld    drain  d1   {Ld*if(dgfs==99,0,1)}

Rth1  Tj      t1              {1.04+limit(Zthtype,0,1)*389.87m}
Rth2  t1      t2              {2.96+limit(Zthtype,0,1)*1.09}
Rth3  t2      t3              {14.09+limit(Zthtype,0,1)*12.96}
Rth4  t3      t4              {73.48+limit(Zthtype,0,1)*47.39}
Rth5  t4      Tcase           {80+limit(Zthtype,0,1)*51.6}
Cth1  Tj      0               3.529u
Cth2  t1      0               1.042u
Cth3  t2      0               1u
Cth4  t3      0               374u
Cth5  t4      0               4.7m


.ENDS
*$



.SUBCKT BSS131_L1 drain gate source PARAMS: dVth=0 dRdson=0 dgfs=0 dC=0

.PARAM Rs=0.074     Rg=10        Ls=3n        Ld=1n        Lg=3n
.PARAM Inn=0.1      Unn=10       Rmax=14
.PARAM act=0.28

X1  d1 g s Tj K_240_a_var PARAMS: a={act} dVth={dVth} dR={dRdson} Inn={Inn} Unn={Unn} 
                                        +Rmax={Rmax} dgfs={dgfs} Rs={Rs} dC={dC} heat=0
Rg    g1     g    {Rg}   
Lg    gate   g1   {Lg*if(dgfs==99,0,1)}
Gs    s1     s    VALUE={V(s1,s)/(Rs*(1+(limit(V(Tj),-200,999)-25)*4m))}
Rsa   s1     s    1Meg
Ls    source s1   {Ls*if(dgfs==99,0,1)}
Ld    drain  d1   {Ld*if(dgfs==99,0,1)}

E1    Tj     w      VALUE={TEMP}
R1    w      0      1u

.ENDS
*$

**********

.SUBCKT BSS87_L1 drain gate source PARAMS: dVth=0 dRdson=0 dgfs=0 dC=0

.PARAM Rs=0.082     Rg=10        Ls=3n        Ld=1n        Lg=3n
.PARAM Inn=0.26     Unn=10       Rmax=6
.PARAM act=0.54

X1  d1 g s Tj K_240_b_var PARAMS: a={act} dVth={dVth} dR={dRdson} Inn={Inn} Unn={Unn} 
                                        +Rmax={Rmax} dgfs={dgfs} Rs={Rs} dC={dC} heat=0
Rg    g1     g    {Rg}   
Lg    gate   g1   {Lg*if(dgfs==99,0,1)}
Gs    s1     s    VALUE={V(s1,s)/(Rs*(1+(limit(V(Tj),-200,999)-25)*4m))}
Rsa   s1     s    1Meg
Ls    source s1   {Ls*if(dgfs==99,0,1)}
Ld    drain  d1   {Ld*if(dgfs==99,0,1)}

E1    Tj     w      VALUE={TEMP}
R1    w      0      1u

.ENDS
*$

**********

.SUBCKT BSP89_L1 drain gate source PARAMS: dVth=0 dRdson=0 dgfs=0 dC=0

.PARAM Rs=0.027     Rg=10        Ls=3n        Ld=1n        Lg=3n
.PARAM Inn=0.35     Unn=10       Rmax=6
.PARAM act=0.54

X1  d1 g s Tj K_240_b_var PARAMS: a={act} dVth={dVth} dR={dRdson} Inn={Inn} Unn={Unn} 
                                        +Rmax={Rmax} dgfs={dgfs} Rs={Rs} dC={dC} heat=0
Rg    g1     g    {Rg}   
Lg    gate   g1   {Lg*if(dgfs==99,0,1)}
Gs    s1     s    VALUE={V(s1,s)/(Rs*(1+(limit(V(Tj),-200,999)-25)*4m))}
Rsa   s1     s    1Meg
Ls    source s1   {Ls*if(dgfs==99,0,1)}
Ld    drain  d1   {Ld*if(dgfs==99,0,1)}

E1    Tj     w      VALUE={TEMP}
R1    w      0      1u

.ENDS
*$

**********

.SUBCKT BSP88_L1 drain gate source PARAMS: dVth=0 dRdson=0 dgfs=0 dC=0

.PARAM Rs=0.027     Rg=10        Ls=3n        Ld=1n        Lg=3n
.PARAM Inn=0.35     Unn=10       Rmax=6
.PARAM act=0.54

X1  d1 g s Tj K_240_c_var PARAMS: a={act} dVth={dVth} dR={dRdson} Inn={Inn} Unn={Unn} 
                                        +Rmax={Rmax} dgfs={dgfs} Rs={Rs} dC={dC} heat=0
Rg    g1     g    {Rg}   
Lg    gate   g1   {Lg*if(dgfs==99,0,1)}
Gs    s1     s    VALUE={V(s1,s)/(Rs*(1+(limit(V(Tj),-200,999)-25)*4m))}
Rsa   s1     s    1Meg
Ls    source s1   {Ls*if(dgfs==99,0,1)}
Ld    drain  d1   {Ld*if(dgfs==99,0,1)}

E1    Tj     w      VALUE={TEMP}
R1    w      0      1u

.ENDS
*$

**********

.SUBCKT BSP129_L1a drain gate source PARAMS: dVth=0 dRdson=0 dgfs=0 dC=0

.PARAM Rs=0.027     Rg=10        Ls=3n        Ld=1n        Lg=3n
.PARAM Inn=0.025    Unn=0        Rmax=20
.PARAM act=0.54

X1  d1 g s Tj K_240_d_var PARAMS: a={act} dVth={dVth} dR={dRdson} Inn={Inn} Unn={Unn} 
                                        +Rmax={Rmax} dgfs={dgfs} Rs={Rs} dC={dC} heat=0
Rg    g1     g    {Rg}   
Lg    gate   g1   {Lg*if(dgfs==99,0,1)}
Gs    s1     s    VALUE={V(s1,s)/(Rs*(1+(limit(V(Tj),-200,999)-25)*4m))}
Rsa   s1     s    1Meg
Ls    source s1   {Ls*if(dgfs==99,0,1)}
Ld    drain  d1   {Ld*if(dgfs==99,0,1)}

E1    Tj     w      VALUE={TEMP}
R1    w      0      1u

.ENDS
*$

**********

.SUBCKT SISC0_97N24D_L1 drain gate source PARAMS: dVth=0 dRdson=0 dgfs=0 dC=0

.PARAM Rs=0.005     Rg=10
.PARAM Inn=0.025    Unn=0        Rmax=20
.PARAM act=0.54

X1  drain g s Tj K_240_d_var PARAMS: a={act} dVth={dVth} dR={dRdson} Inn={Inn} Unn={Unn} 
                                        +Rmax={Rmax} dgfs={dgfs} Rs={Rs} dC={dC} heat=0
Rg    gate     g    {Rg}   

Gs    source     s    VALUE={V(source,s)/(Rs*(1+(limit(V(Tj),-200,999)-25)*4m))}
Rsa   source     s    1Meg

E1    Tj     w      VALUE={TEMP}
R1    w      0      1u

.ENDS

**********

.SUBCKT BSS139_L1 drain gate source PARAMS: dVth=0 dRdson=0 dgfs=0 dC=0

.PARAM Rs=0.074     Rg=10        Ls=3n        Ld=1n        Lg=3n
.PARAM Inn=0.015    Unn=0        Rmax=30
.PARAM act=0.28

X1  d1 g s Tj K_250_d_var PARAMS: a={act} dVth={dVth} dR={dRdson} Inn={Inn} Unn={Unn} 
                                        +Rmax={Rmax} dgfs={dgfs} Rs={Rs} dC={dC} heat=0
Rg    g1     g    {Rg}   
Lg    gate   g1   {Lg*if(dgfs==99,0,1)}
Gs    s1     s    VALUE={V(s1,s)/(Rs*(1+(limit(V(Tj),-200,999)-25)*4m))}
Rsa   s1     s    1Meg
Ls    source s1   {Ls*if(dgfs==99,0,1)}
Ld    drain  d1   {Ld*if(dgfs==99,0,1)}

E1    Tj     w      VALUE={TEMP}
R1    w      0      1u

.ENDS
*$

**********

.SUBCKT BSP324_L1 drain gate source PARAMS: dVth=0 dRdson=0 dgfs=0 dC=0

.PARAM Rs=0.027     Rg=10        Ls=3n        Ld=1n        Lg=3n
.PARAM Inn=0.17     Unn=10       Rmax=25
.PARAM act=0.47

X1  d1 g s Tj K_400_a_var PARAMS: a={act} dVth={dVth} dR={dRdson} Inn={Inn} Unn={Unn} 
                                        +Rmax={Rmax} dgfs={dgfs} Rs={Rs} dC={dC} heat=0
Rg    g1     g    {Rg}   
Lg    gate   g1   {Lg*if(dgfs==99,0,1)}
Gs    s1     s    VALUE={V(s1,s)/(Rs*(1+(limit(V(Tj),-200,999)-25)*4m))}
Rsa   s1     s    1Meg
Ls    source s1   {Ls*if(dgfs==99,0,1)}
Ld    drain  d1   {Ld*if(dgfs==99,0,1)}

E1    Tj     w      VALUE={TEMP}
R1    w      0      1u

.ENDS
*$

**********

.SUBCKT SISC1_4N40E_L1 drain gate source PARAMS: dVth=0 dRdson=0 dgfs=0 dC=0

.PARAM Rs=0.005     Rg=10        
.PARAM Inn=0.17     Unn=10       Rmax=25
.PARAM act=0.47

X1  drain g s Tj K_400_a_var PARAMS: a={act} dVth={dVth} dR={dRdson} Inn={Inn} Unn={Unn} 
                                        +Rmax={Rmax} dgfs={dgfs} Rs={Rs} dC={dC} heat=0
Rg    gate     g    {Rg}   

Gs    source     s    VALUE={V(source,s)/(Rs*(1+(limit(V(Tj),-200,999)-25)*4m))}
Rsa   source     s    1Meg



E1    Tj     w      VALUE={TEMP}
R1    w      0      1u

.ENDS
*$

**********

.SUBCKT BSP125_L1 drain gate source PARAMS: dVth=0 dRdson=0 dgfs=0 dC=0

.PARAM Rs=0.027     Rg=10        Ls=3n        Ld=1n        Lg=3n
.PARAM Inn=0.12     Unn=10       Rmax=45
.PARAM act=0.47

X1  d1 g s Tj K_600_a_var PARAMS: a={act} dVth={dVth} dR={dRdson} Inn={Inn} Unn={Unn} 
                                        +Rmax={Rmax} dgfs={dgfs} Rs={Rs} dC={dC} heat=0
Rg    g1     g    {Rg}   
Lg    gate   g1   {Lg*if(dgfs==99,0,1)}
Gs    s1     s    VALUE={V(s1,s)/(Rs*(1+(limit(V(Tj),-200,999)-25)*4m))}
Rsa   s1     s    1Meg
Ls    source s1   {Ls*if(dgfs==99,0,1)}
Ld    drain  d1   {Ld*if(dgfs==99,0,1)}

E1    Tj     w      VALUE={TEMP}
R1    w      0      1u

.ENDS
*$

**********

.SUBCKT BSS225_L1 drain gate source PARAMS: dVth=0 dRdson=0 dgfs=0 dC=0

.PARAM Rs=0.027     Rg=10        Ls=3n        Ld=1n        Lg=3n
.PARAM Inn=0.12     Unn=10       Rmax=45
.PARAM act=0.47

X1  d1 g s Tj K_600_a_var PARAMS: a={act} dVth={dVth} dR={dRdson} Inn={Inn} Unn={Unn} 
                                        +Rmax={Rmax} dgfs={dgfs} Rs={Rs} dC={dC} heat=0
Rg    g1     g    {Rg}   
Lg    gate   g1   {Lg*if(dgfs==99,0,1)}
Gs    s1     s    VALUE={V(s1,s)/(Rs*(1+(limit(V(Tj),-200,999)-25)*4m))}
Rsa   s1     s    1Meg
Ls    source s1   {Ls*if(dgfs==99,0,1)}
Ld    drain  d1   {Ld*if(dgfs==99,0,1)}

E1    Tj     w      VALUE={TEMP}
R1    w      0      1u

.ENDS

**********

.SUBCKT BSS127_L1 drain gate source PARAMS: dVth=0 dRdson=0 dgfs=0 dC=0

.PARAM Rs=0.074     Rg=10        Ls=3n        Ld=1n        Lg=3n
.PARAM Inn=0.016    Unn=10       Rmax=500
.PARAM act=0.04

X1  d1 g s Tj K_600_a_var PARAMS: a={act} dVth={dVth} dR={dRdson} Inn={Inn} Unn={Unn} 
                                        +Rmax={Rmax} dgfs={dgfs} Rs={Rs} dC={dC} heat=0
Rg    g1     g    {Rg}   
Lg    gate   g1   {Lg*if(dgfs==99,0,1)}
Gs    s1     s    VALUE={V(s1,s)/(Rs*(1+(limit(V(Tj),-200,999)-25)*4m))}
Rsa   s1     s    1Meg
Ls    source s1   {Ls*if(dgfs==99,0,1)}
Ld    drain  d1   {Ld*if(dgfs==99,0,1)}

E1    Tj     w      VALUE={TEMP}
R1    w      0      1u

.ENDS

**********

.SUBCKT BSP135_L1 drain gate source PARAMS: dVth=0 dRdson=0 dgfs=0 dC=0

.PARAM Rs=0.027     Rg=10        Ls=3n        Ld=1n        Lg=3n
.PARAM Inn=0.01     Unn=0        Rmax=60
.PARAM act=0.47

X1  d1 g s Tj K_600_d_var PARAMS: a={act} dVth={dVth} dR={dRdson} Inn={Inn} Unn={Unn} 
                                        +Rmax={Rmax} dgfs={dgfs} Rs={Rs} dC={dC} heat=0
Rg    g1     g    {Rg}   
Lg    gate   g1   {Lg*if(dgfs==99,0,1)}
Gs    s1     s    VALUE={V(s1,s)/(Rs*(1+(limit(V(Tj),-200,999)-25)*4m))}
Rsa   s1     s    1Meg
Ls    source s1   {Ls*if(dgfs==99,0,1)}
Ld    drain  d1   {Ld*if(dgfs==99,0,1)}

E1    Tj     w      VALUE={TEMP}
R1    w      0      1u

.ENDS
*$

**********

.SUBCKT SISC1_4N60D_L1 drain gate source PARAMS: dVth=0 dRdson=0 dgfs=0 dC=0

.PARAM Rs=0.005     Rg=10        
.PARAM Inn=0.01     Unn=0        Rmax=60
.PARAM act=0.47

X1  drain g s Tj K_600_d_var PARAMS: a={act} dVth={dVth} dR={dRdson} Inn={Inn} Unn={Unn} 
                                        +Rmax={Rmax} dgfs={dgfs} Rs={Rs} dC={dC} heat=0
Rg    gate     g    {Rg}   

Gs    source     s    VALUE={V(source,s)/(Rs*(1+(limit(V(Tj),-200,999)-25)*4m))}
Rsa   source     s    1Meg



E1    Tj     w      VALUE={TEMP}
R1    w      0      1u

.ENDS

**********

.SUBCKT BSS126_L1 drain gate source PARAMS: dVth=0 dRdson=0 dgfs=0 dC=0

.PARAM Rs=0.074     Rg=0.9       Ls=3n        Ld=1n        Lg=3n
.PARAM Inn=0.003    Unn=0        Rmax=700
.PARAM act=0.04

X1  d1 g s Tj K_600_e_var PARAMS: a={act} dVth={dVth} dR={dRdson} Inn={Inn} Unn={Unn} 
                                        +Rmax={Rmax} dgfs={dgfs} Rs={Rs} dC={dC} heat=0
Rg    g1     g    {Rg}   
Lg    gate   g1   {Lg*if(dgfs==99,0,1)}
Gs    s1     s    VALUE={V(s1,s)/(Rs*(1+(limit(V(Tj),-200,999)-25)*4m))}
Rsa   s1     s    1Meg
Ls    source s1   {Ls*if(dgfs==99,0,1)}
Ld    drain  d1   {Ld*if(dgfs==99,0,1)}

E1    Tj     w      VALUE={TEMP}
R1    w      0      1u

.ENDS

**********

.SUBCKT BSS131_L0  drain  gate  source

Lg     gate  g1    3n
Ld     drain d1    1n
Ls     source s1   3n
Rs      s1    s2   0.074

Rg     g1    g2     10
M1      d2    g2    s2    s2    DMOS    L=1u   W=1u
.MODEL DMOS NMOS ( KP= 0.223  VTO=1.6  THETA=0  VMAX=1.5e5  ETA=0  LEVEL=3)
Rd     d2    d1a    6.07 TC=11m
.MODEL MVDR NMOS (KP=0.55 VTO=-1.4   LAMBDA=0.15)
Mr d1 d2a d1a d1a MVDR W=1u L=1u
Rx d2a d1a 1m

Dbd     s2    d2    Dbt
.MODEL     Dbt    D(BV=290   M=0.5  CJO=34.44p  VJ=0.5V)
Dbody   s2   21    DBODY
.MODEL DBODY  D(IS=7p  N=1.2  RS=475u  EG=1.12  TT=60n)
Rdiode  d1  21    714.29m TC=1m

.MODEL   sw    NMOS(VTO=0  KP=10   LEVEL=1)
Maux      g2   c    a    a   sw
Maux2     b    d    g2    g2   sw
Eaux      c    a    d2    g2   1
Eaux2     d    g2   d2    g2   -1
Cox       b    d2   99.4p
.MODEL     DGD    D(M=1   CJO=99.4p   VJ=0.5)
Rpar      b    d2   1Meg
Dgd       a    d2   DGD
Rpar2     d2   a    10Meg
Cgs     g2    s2    55.44p

.ENDS  BSS131_L0

******

.SUBCKT BSS87_L0  drain  gate  source

Lg     gate  g1    3n
Ld     drain d1    1n
Ls     source s1   3n
Rs      s1    s2   0.082

Rg     g1    g2     10
M1      d2    g2    s2    s2    DMOS    L=1u   W=1u
.MODEL DMOS NMOS ( KP= 0.486  VTO=1.7  THETA=0  VMAX=1.5e5  ETA=0  LEVEL=3)
Rd     d2    d1a    3.15 TC=11m
.MODEL MVDR NMOS (KP=1.05 VTO=-1.4   LAMBDA=0.15)
Mr d1 d2a d1a d1a MVDR W=1u L=1u
Rx d2a d1a 1m

Dbd     s2    d2    Dbt
.MODEL     Dbt    D(BV=290   M=0.5  CJO=66.42p  VJ=0.5V)
Dbody   s2   21    DBODY
.MODEL DBODY  D(IS=13.5p  N=1.2  RS=246u  EG=1.12  TT=60n)
Rdiode  d1  21    370.37m TC=1m

.MODEL   sw    NMOS(VTO=0  KP=10   LEVEL=1)
Maux      g2   c    a    a   sw
Maux2     b    d    g2    g2   sw
Eaux      c    a    d2    g2   1
Eaux2     d    g2   d2    g2   -1
Cox       b    d2   180.9p
.MODEL     DGD    D(M=0.76   CJO=180.9p   VJ=0.5)
Rpar      b    d2   1Meg
Dgd       a    d2   DGD
Rpar2     d2   a    10Meg
Cgs     g2    s2    75.06p

.ENDS  BSS87_L0

******

.SUBCKT BSP89_L0  drain  gate  source

Lg     gate  g1    3n
Ld     drain d1    1n
Ls     source s1   3n
Rs      s1    s2   0.027

Rg     g1    g2     10
M1      d2    g2    s2    s2    DMOS    L=1u   W=1u
.MODEL DMOS NMOS ( KP= 0.486  VTO=1.7  THETA=0  VMAX=1.5e5  ETA=0  LEVEL=3)
Rd     d2    d1a    3.15 TC=11m
.MODEL MVDR NMOS (KP=1.05 VTO=-1.4   LAMBDA=0.15)
Mr d1 d2a d1a d1a MVDR W=1u L=1u
Rx d2a d1a 1m

Dbd     s2    d2    Dbt
.MODEL     Dbt    D(BV=290   M=0.5  CJO=66.42p  VJ=0.5V)
Dbody   s2   21    DBODY
.MODEL DBODY  D(IS=13.5p  N=1.2  RS=246u  EG=1.12  TT=60n)
Rdiode  d1  21    370.37m TC=1m

.MODEL   sw    NMOS(VTO=0  KP=10   LEVEL=1)
Maux      g2   c    a    a   sw
Maux2     b    d    g2    g2   sw
Eaux      c    a    d2    g2   1
Eaux2     d    g2   d2    g2   -1
Cox       b    d2   180.9p
.MODEL     DGD    D(M=0.76   CJO=180.9p   VJ=0.5)
Rpar      b    d2   1Meg
Dgd       a    d2   DGD
Rpar2     d2   a    10Meg
Cgs     g2    s2    75.06p

.ENDS  BSP89_L0

******

.SUBCKT BSP88_L0  drain  gate  source

Lg     gate  g1    3n
Ld     drain d1    1n
Ls     source s1   3n
Rs      s1    s2   0.027

Rg     g1    g2     10
M1      d2    g2    s2    s2    DMOS    L=1u   W=1u
.MODEL DMOS NMOS ( KP= 0.486  VTO=1.3  THETA=0  VMAX=1.5e5  ETA=0  LEVEL=3)
Rd     d2    d1a    3.15 TC=11m
.MODEL MVDR NMOS (KP=0.89 VTO=-1.4   LAMBDA=0.15)
Mr d1 d2a d1a d1a MVDR W=1u L=1u
Rx d2a d1a 1m

Dbd     s2    d2    Dbt
.MODEL     Dbt    D(BV=290   M=0.5  CJO=66.42p  VJ=0.5V)
Dbody   s2   21    DBODY
.MODEL DBODY  D(IS=13.5p  N=1.2  RS=246u  EG=1.12  TT=60n)
Rdiode  d1  21    370.37m TC=1m

.MODEL   sw    NMOS(VTO=0  KP=10   LEVEL=1)
Maux      g2   c    a    a   sw
Maux2     b    d    g2    g2   sw
Eaux      c    a    d2    g2   1
Eaux2     d    g2   d2    g2   -1
Cox       b    d2   180.9p
.MODEL     DGD    D(M=0.77   CJO=180.9p   VJ=0.5)
Rpar      b    d2   1Meg
Dgd       a    d2   DGD
Rpar2     d2   a    10Meg
Cgs     g2    s2    75.06p

.ENDS  BSP88_L0

******

.SUBCKT BSP129_L0  drain  gate  source

Lg     gate  g1    3n
Ld     drain d1    1n
Ls     source s1   3n
Rs      s1    s2   0.027

Rg     g1    g2     10
M1      d2    g2    s2    s2    DMOS    L=1u   W=1u
.MODEL DMOS NMOS ( KP= 0.486  VTO=-0.85  THETA=0  VMAX=1.5e5  ETA=0  LEVEL=3)
Rd     d2    d1a    3.15 TC=11m
.MODEL MVDR NMOS (KP=1.05 VTO=-1.4   LAMBDA=0.15)
Mr d1 d2a d1a d1a MVDR W=1u L=1u
Rx d2a d1a 1m

Dbd     s2    d2    Dbt
.MODEL     Dbt    D(BV=290   M=0.5  CJO=66.42p  VJ=0.5V)
Dbody   s2   21    DBODY
.MODEL DBODY  D(IS=13.5p  N=1.2  RS=246u  EG=1.12  TT=60n)
Rdiode  d1  21    370.37m TC=1m

.MODEL   sw    NMOS(VTO=0  KP=10   LEVEL=1)
Maux      g2   c    a    a   sw
Maux2     b    d    g2    g2   sw
Eaux      c    a    d2    g2   1
Eaux2     d    g2   d2    g2   -1
Cox       b    d2   180.9p
.MODEL     DGD    D(M=0.66   CJO=180.9p   VJ=0.5)
Rpar      b    d2   1Meg
Dgd       a    d2   DGD
Rpar2     d2   a    10Meg
Cgs     g2    s2    75.06p

.ENDS  BSP129_L0

******

.SUBCKT SISC0_97N24D_L0  drain  gate  source




Rs      source    s2   0.005

Rg     gate    g2     10
M1      d2    g2    s2    s2    DMOS    L=1u   W=1u
.MODEL DMOS NMOS ( KP= 0.486  VTO=-0.85  THETA=0  VMAX=1.5e5  ETA=0  LEVEL=3)
Rd     d2    d1a    3.15 TC=11m
.MODEL MVDR NMOS (KP=1.05 VTO=-1.4   LAMBDA=0.15)
Mr drain d2a d1a d1a MVDR W=1u L=1u
Rx d2a d1a 1m

Dbd     s2    d2    Dbt
.MODEL     Dbt    D(BV=290   M=0.5  CJO=66.42p  VJ=0.5V)
Dbody   s2   21    DBODY
.MODEL DBODY  D(IS=13.5p  N=1.2  RS=246u  EG=1.12  TT=60n)
Rdiode  drain  21    370.37m TC=1m

.MODEL   sw    NMOS(VTO=0  KP=10   LEVEL=1)
Maux      g2   c    a    a   sw
Maux2     b    d    g2    g2   sw
Eaux      c    a    d2    g2   1
Eaux2     d    g2   d2    g2   -1
Cox       b    d2   180.9p
.MODEL     DGD    D(M=0.66   CJO=180.9p   VJ=0.5)
Rpar      b    d2   1Meg
Dgd       a    d2   DGD
Rpar2     d2   a    10Meg
Cgs     g2    s2    75.06p

.ENDS  SISC0_97N24D_L0

******

.SUBCKT BSS139_L0  drain  gate  source

Lg     gate  g1    3n
Ld     drain d1    1n
Ls     source s1   3n
Rs      s1    s2   0.074

Rg     g1    g2     10
M1      d2    g2    s2    s2    DMOS    L=1u   W=1u
.MODEL DMOS NMOS ( KP= 0.223  VTO=-0.89  THETA=0  VMAX=1.5e5  ETA=0  LEVEL=3)
Rd     d2    d1a    7.14 TC=11m
.MODEL MVDR NMOS (KP=0.55 VTO=-1.4   LAMBDA=0.15)
Mr d1 d2a d1a d1a MVDR W=1u L=1u
Rx d2a d1a 1m

Dbd     s2    d2    Dbt
.MODEL     Dbt    D(BV=295   M=0.5  CJO=34.44p  VJ=0.5V)
Dbody   s2   21    DBODY
.MODEL DBODY  D(IS=7p  N=1.2  RS=475u  EG=1.12  TT=60n)
Rdiode  d1  21    714.29m TC=1m

.MODEL   sw    NMOS(VTO=0  KP=10   LEVEL=1)
Maux      g2   c    a    a   sw
Maux2     b    d    g2    g2   sw
Eaux      c    a    d2    g2   1
Eaux2     d    g2   d2    g2   -1
Cox       b    d2   106.12p
.MODEL     DGD    D(M=0.66   CJO=106.12p   VJ=0.5)
Rpar      b    d2   1Meg
Dgd       a    d2   DGD
Rpar2     d2   a    10Meg
Cgs     g2    s2    55.44p

.ENDS  BSS139_L0

******

.SUBCKT BSP324_L0  drain  gate  source

Lg     gate  g1    3n
Ld     drain d1    1n
Ls     source s1   3n
Rs      s1    s2   0.027

Rg     g1    g2     10
M1      d2    g2    s2    s2    DMOS    L=1u   W=1u
.MODEL DMOS NMOS ( KP= 0.273  VTO=2.27  THETA=0  VMAX=1.5e5  ETA=0  LEVEL=3)
Rd     d2    d1a    12.23 TC=11m
.MODEL MVDR NMOS (KP=0.4 VTO=-1.4   LAMBDA=0.15)
Mr d1 d2a d1a d1a MVDR W=1u L=1u
Rx d2a d1a 1m

Dbd     s2    d2    Dbt
.MODEL     Dbt    D(BV=495   M=0.5  CJO=57.81p  VJ=0.5V)
Dbody   s2   21    DBODY
.MODEL DBODY  D(IS=11.8p  N=1.2  RS=283u  EG=1.12  TT=80n)
Rdiode  d1  21    425.53m TC=0

.MODEL   sw    NMOS(VTO=0  KP=10   LEVEL=1)
Maux      g2   c    a    a   sw
Maux2     b    d    g2    g2   sw
Eaux      c    a    d2    g2   1
Eaux2     d    g2   d2    g2   -1
Cox       b    d2   220.9p
.MODEL     DGD    D(M=0.97   CJO=220.9p   VJ=0.5)
Rpar      b    d2   1Meg
Dgd       a    d2   DGD
Rpar2     d2   a    10Meg
Cgs     g2    s2    95.88p

.ENDS  BSP324_L0

******

.SUBCKT SISC1_4N40E_L0  drain  gate  source




Rs      source    s2   0.005

Rg     gate    g2     10
M1      d2    g2    s2    s2    DMOS    L=1u   W=1u
.MODEL DMOS NMOS ( KP= 0.273  VTO=2.27  THETA=0  VMAX=1.5e5  ETA=0  LEVEL=3)
Rd     d2    d1a    12.23 TC=11m
.MODEL MVDR NMOS (KP=0.4 VTO=-1.4   LAMBDA=0.15)
Mr drain d2a d1a d1a MVDR W=1u L=1u
Rx d2a d1a 1m

Dbd     s2    d2    Dbt
.MODEL     Dbt    D(BV=495   M=0.5  CJO=57.81p  VJ=0.5V)
Dbody   s2   21    DBODY
.MODEL DBODY  D(IS=11.8p  N=1.2  RS=283u  EG=1.12  TT=80n)
Rdiode  drain  21    425.53m TC=0

.MODEL   sw    NMOS(VTO=0  KP=10   LEVEL=1)
Maux      g2   c    a    a   sw
Maux2     b    d    g2    g2   sw
Eaux      c    a    d2    g2   1
Eaux2     d    g2   d2    g2   -1
Cox       b    d2   220.9p
.MODEL     DGD    D(M=0.97   CJO=220.9p   VJ=0.5)
Rpar      b    d2   1Meg
Dgd       a    d2   DGD
Rpar2     d2   a    10Meg
Cgs     g2    s2    95.88p

.ENDS  SISC1_4N40E_L0

******

.SUBCKT BSP125_L0  drain  gate  source

Lg     gate  g1    3n
Ld     drain d1    1n
Ls     source s1   3n
Rs      s1    s2   0.027

Rg     g1    g2     10
M1      d2    g2    s2    s2    DMOS    L=1u   W=1u
.MODEL DMOS NMOS ( KP= 0.273  VTO=2.27  THETA=0  VMAX=1.5e5  ETA=0  LEVEL=3)
Rd     d2    d1a    23.4 TC=11m
.MODEL MVDR NMOS (KP=0.24 VTO=-1.4   LAMBDA=0.15)
Mr d1 d2a d1a d1a MVDR W=1u L=1u
Rx d2a d1a 1m

Dbd     s2    d2    Dbt
.MODEL     Dbt    D(BV=650   M=0.5  CJO=57.81p  VJ=0.5V)
Dbody   s2   21    DBODY
.MODEL DBODY  D(IS=11.8p  N=1.2  RS=283u  EG=1.12  TT=130n)
Rdiode  d1  21    425.53m TC=0

.MODEL   sw    NMOS(VTO=0  KP=10   LEVEL=1)
Maux      g2   c    a    a   sw
Maux2     b    d    g2    g2   sw
Eaux      c    a    d2    g2   1
Eaux2     d    g2   d2    g2   -1
Cox       b    d2   220.9p
.MODEL     DGD    D(M=1   CJO=220.9p   VJ=0.5)
Rpar      b    d2   1Meg
Dgd       a    d2   DGD
Rpar2     d2   a    10Meg
Cgs     g2    s2    95.88p

.ENDS  BSP125_L0

******

.SUBCKT BSS225_L0  drain  gate  source

Lg     gate  g1    3n
Ld     drain d1    1n
Ls     source s1   3n
Rs      s1    s2   0.027

Rg     g1    g2     10
M1      d2    g2    s2    s2    DMOS    L=1u   W=1u
.MODEL DMOS NMOS ( KP= 0.273  VTO=2.27  THETA=0  VMAX=1.5e5  ETA=0  LEVEL=3)
Rd     d2    d1a    23.4 TC=11m
.MODEL MVDR NMOS (KP=0.24 VTO=-1.4   LAMBDA=0.15)
Mr d1 d2a d1a d1a MVDR W=1u L=1u
Rx d2a d1a 1m

Dbd     s2    d2    Dbt
.MODEL     Dbt    D(BV=650   M=0.5  CJO=57.81p  VJ=0.5V)
Dbody   s2   21    DBODY
.MODEL DBODY  D(IS=11.8p  N=1.2  RS=283u  EG=1.12  TT=130n)
Rdiode  d1  21    425.53m TC=0

.MODEL   sw    NMOS(VTO=0  KP=10   LEVEL=1)
Maux      g2   c    a    a   sw
Maux2     b    d    g2    g2   sw
Eaux      c    a    d2    g2   1
Eaux2     d    g2   d2    g2   -1
Cox       b    d2   220.9p
.MODEL     DGD    D(M=1   CJO=220.9p   VJ=0.5)
Rpar      b    d2   1Meg
Dgd       a    d2   DGD
Rpar2     d2   a    10Meg
Cgs     g2    s2    95.88p

.ENDS  BSS225_L0

******

.SUBCKT BSP135_L0  drain  gate  source

Lg     gate  g1    3n
Ld     drain d1    1n
Ls     source s1   3n
Rs      s1    s2   0.027

Rg     g1    g2     10
M1      d2    g2    s2    s2    DMOS    L=1u   W=1u
.MODEL DMOS NMOS ( KP= 0.273  VTO=-0.93  THETA=0  VMAX=1.5e5  ETA=0  LEVEL=3)
Rd     d2    d1a    21.91 TC=11m
.MODEL MVDR NMOS (KP=0.24 VTO=-1.4   LAMBDA=0.15)
Mr d1 d2a d1a d1a MVDR W=1u L=1u
Rx d2a d1a 1m

Dbd     s2    d2    Dbt
.MODEL     Dbt    D(BV=650   M=0.5  CJO=57.81p  VJ=0.5V)
Dbody   s2   21    DBODY
.MODEL DBODY  D(IS=11.8p  N=1.2  RS=283u  EG=1.12  TT=130n)
Rdiode  d1  21    425.53m TC=0

.MODEL   sw    NMOS(VTO=0  KP=10   LEVEL=1)
Maux      g2   c    a    a   sw
Maux2     b    d    g2    g2   sw
Eaux      c    a    d2    g2   1
Eaux2     d    g2   d2    g2   -1
Cox       b    d2   213.85p
.MODEL     DGD    D(M=0.7   CJO=213.85p   VJ=0.5)
Rpar      b    d2   1Meg
Dgd       a    d2   DGD
Rpar2     d2   a    10Meg
Cgs     g2    s2    95.88p

.ENDS  BSP135_L0

******

.SUBCKT SISC1_4N60D_L0  drain  gate  source




Rs      source    s2   0.005

Rg     gate    g2     10
M1      d2    g2    s2    s2    DMOS    L=1u   W=1u
.MODEL DMOS NMOS ( KP= 0.273  VTO=-0.93  THETA=0  VMAX=1.5e5  ETA=0  LEVEL=3)
Rd     d2    d1a    21.91 TC=11m
.MODEL MVDR NMOS (KP=0.24 VTO=-1.4   LAMBDA=0.15)
Mr drain d2a d1a d1a MVDR W=1u L=1u
Rx d2a d1a 1m

Dbd     s2    d2    Dbt
.MODEL     Dbt    D(BV=650   M=0.5  CJO=57.81p  VJ=0.5V)
Dbody   s2   21    DBODY
.MODEL DBODY  D(IS=11.8p  N=1.2  RS=283u  EG=1.12  TT=130n)
Rdiode  drain  21    425.53m TC=0

.MODEL   sw    NMOS(VTO=0  KP=10   LEVEL=1)
Maux      g2   c    a    a   sw
Maux2     b    d    g2    g2   sw
Eaux      c    a    d2    g2   1
Eaux2     d    g2   d2    g2   -1
Cox       b    d2   213.85p
.MODEL     DGD    D(M=0.7   CJO=213.85p   VJ=0.5)
Rpar      b    d2   1Meg
Dgd       a    d2   DGD
Rpar2     d2   a    10Meg
Cgs     g2    s2    95.88p

.ENDS  SISC1_4N60D_L0

******

.SUBCKT BSS127_L0  drain  gate  source

Lg     gate  g1    3n
Ld     drain d1    1n
Ls     source s1   3n
Rs      s1    s2   0.074

Rg     g1    g2     10
M1      d2    g2    s2    s2    DMOS    L=1u   W=1u
.MODEL DMOS NMOS ( KP= 0.023  VTO=2.27  THETA=0  VMAX=1.5e5  ETA=0  LEVEL=3)
Rd     d2    d1a    275 TC=11m
.MODEL MVDR NMOS (KP=0.02 VTO=-1.4   LAMBDA=0.15)
Mr d1 d2a d1a d1a MVDR W=1u L=1u
Rx d2a d1a 1m

Dbd     s2    d2    Dbt
.MODEL     Dbt    D(BV=650   M=0.5  CJO=4.92p  VJ=0.5V)
Dbody   s2   21    DBODY
.MODEL DBODY  D(IS=1p  N=1.2  RS=3325u  EG=1.12  TT=130n)
Rdiode  d1  21    5000m TC=0

.MODEL   sw    NMOS(VTO=0  KP=10   LEVEL=1)
Maux      g2   c    a    a   sw
Maux2     b    d    g2    g2   sw
Eaux      c    a    d2    g2   1
Eaux2     d    g2   d2    g2   -1
Cox       b    d2   18.8p
.MODEL     DGD    D(M=1   CJO=18.8p   VJ=0.5)
Rpar      b    d2   1Meg
Dgd       a    d2   DGD
Rpar2     d2   a    10Meg
Cgs     g2    s2    8.16p

.ENDS  BSS127_L0

******

.SUBCKT BSS126_L0  drain  gate  source

Lg     gate  g1    3n
Ld     drain d1    1n
Ls     source s1   3n
Rs      s1    s2   0.074

Rg     g1    g2     10
M1      d2    g2    s2    s2    DMOS    L=1u   W=1u
.MODEL DMOS NMOS ( KP= 0.03  VTO=-1.53  THETA=0  VMAX=1.5e5  ETA=0  LEVEL=3)
Rd     d2    d1a    275 TC=11m
.MODEL MVDR NMOS (KP=0.02 VTO=-1.4   LAMBDA=0.15)
Mr d1 d2a d1a d1a MVDR W=1u L=1u
Rx d2a d1a 1m

Dbd     s2    d2    Dbt
.MODEL     Dbt    D(BV=650   M=0.5  CJO=4.92p  VJ=0.5V)
Dbody   s2   21    DBODY
.MODEL DBODY  D(IS=1p  N=1.2  RS=3325u  EG=1.12  TT=130n)
Rdiode  d1  21    5000m TC=0

.MODEL   sw    NMOS(VTO=0  KP=10   LEVEL=1)
Maux      g2   c    a    a   sw
Maux2     b    d    g2    g2   sw
Eaux      c    a    d2    g2   1
Eaux2     d    g2   d2    g2   -1
Cox       b    d2   24p
.MODEL     DGD    D(M=0.6   CJO=24p   VJ=0.5)
Rpar      b    d2   1Meg
Dgd       a    d2   DGD
Rpar2     d2   a    10Meg
Cgs     g2    s2    20p

.ENDS  BSS126_L0

************

.SUBCKT BSP300_L0  drain  gate  source

Lg     gate  g1    3n
Ld     drain d1    2n
Ls     source s1   3n
Rs      s1    s2   0.074

Rg     g1    g2     10
M1      d2    g2    s2    s2    DMOS    L=1u   W=1u
.MODEL DMOS NMOS ( KP= 0.4  VTO=3.4  THETA=0  VMAX=1.5e5  ETA=0  LEVEL=3)
Rd     d2    d1a    15 TC=5.5m

.MODEL MVDR NMOS (KP=3.83 VTO=-1.4   LAMBDA=0.15)
Mr d1 d2a d1a d1a MVDR W=1u L=1u
Rx d2a d1a 1m

Dbd     s2    d2    Dbt
.MODEL     Dbt    D(BV=800   M=0.5  CJO=200p  VJ=0.5V)
Dbody   s2   21    DBODY
.MODEL DBODY  D(IS=3p  N=1  RS=30u  EG=1.12  TT=700n)
Rdiode  d1  21    0.8 TC=0

.MODEL   sw    NMOS(VTO=0  KP=10   LEVEL=1)
Maux      g2   c    a    a   sw
Maux2     b    d    g2    g2   sw
Eaux      c    a    d2    g2   1
Eaux2     d    g2   d2    g2   -1
Cox       b    d2   900p
.MODEL     DGD    D(M=0.97   CJO=400p   VJ=0.5)
Rpar      b    d2   1Meg
Dgd       a    d2   DGD
Rpar2     d2   a    10Meg
Cgs     g2    s2    170p

.ENDS  BSP300_L0

******






**** Netlist ****
Vbat  vb gnd DC 3.9
Vcs   vb col DC 0
Vbias vb bias DC 0
X1    col base gnd KSC5502D 
X2    bias en base BSP125_L0

Ven en gnd DC 0 PWL(0s 0v 0.0004s 0v 0.0007s 3.9v 3s 3.9v) r=0


**** Simulation ****
.tran 0.01m 0.0012s
.control
run
set color0 = white ; plot window - background color
set color1 = black ; plot window - grid and text color
plot I(Vcs) I(Vbias)
plot V(en,base)
print I(Vcs) I(Vbias)
.endc
.end
