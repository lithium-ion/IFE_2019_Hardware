RC Circuit Transient Response
**** Models ****

*---------------------------------------------------------------*
* Panasonic JS-M Automotive SPDT Relay Model
*    
*    Simulate the behavior of the SPDT Relay
*    Caution - No 10ms Delay
*
*                   Positive Side of Coil
*                   |     Negative Side of Coil
*                   |     |      Common
*                   |     |      |     Normally Open
*                   |     |      |     |   Normally Closed
*---------------------------------------------------------------*
.SUBCKT RELAY_SPDT wcoila wcoilb wcom wno wnc
Rcoil wcoila 1 225
Lcoil 1 wcoilb 1uH
S1 wnc wcom wcoila wcoilb swclosed OFF
S2 wcom wno wcoila wcoilb swopen OFF
.model swopen SW vt = 6.3 vh = 5.4 ron = 0.1u roff = 10g
.model swclosed SW vt = 6.3 vh = 5.4 ron = 10g roff = 0.1u
.ends RELAY_SPDT


*---------------------------------------------------------------*
* TE EV200 Contactor Model
*    
*    Simulate the Inrush Current + Steady State Current
*
*                         Positive Side of Coil
*                         |     Negative Side of Coil
*                         |     |
*---------------------------------------------------------------*
.SUBCKT EV200_CONTACTOR coila coilb
Rsteady coila a 123
Lsteady a coilb 100u
.ends EV200_CONTACTOR


*---------------------------------------------------------------*
* LM393 VOLTAGE COMPARATOR "MACROMODEL" SUBCIRCUIT
* CREATED USING PARTS VERSION 4.03 ON 03/07/90 AT 14:17
* REV (N/A)
* CONNECTIONS:   NON-INVERTING INPUT
*                | INVERTING INPUT
*                | | POSITIVE POWER SUPPLY
*                | | | NEGATIVE POWER SUPPLY
*                | | | | OPEN COLLECTOR OUTPUT
*                | | | | |
*---------------------------------------------------------------*
.SUBCKT LM393    1 2 3 4 5
  F1    9  3 V1 1
  IEE   3  7 DC 100.0E-6
  VI1  21  1 DC .75
  VI2  22  2 DC .75
  Q1    9 21  7 QIN
  Q2    8 22  7 QIN
  Q3    9  8  4 QMO
  Q4    8  8  4 QMI
.MODEL QIN PNP(IS=800.0E-18 BF=2.000E3)
.MODEL QMI NPN(IS=800.0E-18 BF=1002)
.MODEL QMO NPN(IS=800.0E-18 BF=1000 CJC=1E-15 TR=807.4E-9)
  E1   10  4  9  4  1
  V1   10 11 DC 0
  Q5    5 11  4 QOC
.MODEL QOC NPN(IS=800.0E-18 BF=20.29E3 CJC=1E-15 TF=942.6E-12 TR=543.8E-9)
  DP    4  3 DX
  RP 3  4 46.3E3
.MODEL DX  D(IS=800.0E-18)
.ENDS LM393



.SUBCKT ntd20n03l27 1 2 3
**************************************
*      Model Generated by MODPEX     *
*Copyright(c) Symmetry Design Systems*
*         All Rights Reserved        *
*    UNPUBLISHED LICENSED SOFTWARE   *
*   Contains Proprietary Information *
*      Which is The Property of      *
*     SYMMETRY OR ITS LICENSORS      *
*Commercial Use or Resale Restricted *
*   by Symmetry License Agreement    *
**************************************
* Model generated on Dec  7, 04
* MODEL FORMAT: PSpice
* Symmetry POWER MOS Model (Version 1.0)
* External Node Designations
* Node 1 -> Drain
* Node 2 -> Gate
* Node 3 -> Source
M1 9 7 8 8 MM L=100u W=100u
* Default values used in MM:
* The voltage-dependent capacitances are
* not included. Other default values are:
*   RS=0 RD=0 LD=0 CBD=0 CBS=0 CGBO=0
.MODEL MM NMOS LEVEL=1 IS=1e-32
+VTO=2.22412 LAMBDA=0.0386082 KP=85.4982
+CGSO=8.95186e-06 CGDO=8.51054e-09
RS 8 3 0.0174624
D1 3 1 MD
.MODEL MD D IS=1e-07 RS=0.00439529 N=1.68776 BV=30
+IBV=0.00025 EG=1.2 XTI=4 TT=0
+CJO=9.31194e-10 VJ=0.499875 M=0.364891 FC=0.5
RDS 3 1 2.77e+11
RD 9 1 0.0001
RG 2 7 18.429
D2 4 5 MD1
* Default values used in MD1:
*   RS=0 EG=1.11 XTI=3.0 TT=0
*   BV=infinite IBV=1mA
.MODEL MD1 D IS=1e-32 N=50
+CJO=6.36264e-10 VJ=1.13275 M=0.76851 FC=9.99812e-09
D3 0 5 MD2
* Default values used in MD2:
*   EG=1.11 XTI=3.0 TT=0 CJO=0
*   BV=infinite IBV=1mA
.MODEL MD2 D IS=1e-10 N=1.39383 RS=2.75597e-06
RL 5 10 1
FI2 7 9 VFI2 -1
VFI2 4 0 0
EV16 10 0 9 7 1
CAP 11 10 6.36264e-10
FI1 7 9 VFI1 -1
VFI1 11 6 0
RCAP 6 10 1
D4 0 6 MD3
* Default values used in MD3:
*   EG=1.11 XTI=3.0 TT=0 CJO=0
*   RS=0 BV=infinite IBV=1mA
.MODEL MD3 D IS=1e-10 N=1.39383
.ENDS ntd20n03l27



**** Netlist ****
Rset vdd n2 7k
Rdist n3 gnd 100
Ru vdd n4 3.7k
Rl n4 gnd 6.3k
R0 vdd gnd 10k
R1 vdd pc_comp 10k
C0 n1 gnd 1000u
X0 vdd gnd n1 n2 n3 RELAY_SPDT
X1 n1 n4 vdd gnd pc_comp LM393
vin vdd gnd DC 0 PULSE(0v 16v 1s 1us 1us 10s) PULSE(0v 16v 10.5s 1us 1us 10s)

X2 vdd n7 EV200_CONTACTOR
Dflyback vdd n7 Da1N4004
.model Da1N4004 D (IS=18.8n RS=0 BV=400 IBV=5.00u CJO=30 M=0.333 N=2)
X3 n7 pc_comp n8 ntd20n03l27
Vdummy n8 gnd 0


**** Simulation ****
.tran 0.1m 15s
.control
run
set color0 = white ; plot window - background color
set color1 = black ; plot window - grid and text color
plot v(vdd) v(n1) v(n4) v(pc_comp)
plot v(pc_comp) v(n7)
.endc
.end
